
library ieee; 
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package Sigmoid_Package is
    TYPE sigmoid_array IS ARRAY (0 to 65535) OF NATURAL range 0 to 65535;
    CONSTANT sigmoid : sigmoid_array := (0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 11, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 12, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 13, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 14, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 16, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 17, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 19, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 20, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 22, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 23, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 25, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 26, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 29, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 51, 51, 51, 51, 51, 51, 51, 51, 51, 51, 51, 51, 51, 51, 51, 51, 51, 51, 51, 51, 51, 51, 51, 51, 51, 51, 51, 51, 51, 51, 51, 51, 51, 51, 51, 51, 51, 51, 51, 51, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 52, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 53, 54, 54, 54, 54, 54, 54, 54, 54, 54, 54, 54, 54, 54, 54, 54, 54, 54, 54, 54, 54, 54, 54, 54, 54, 54, 54, 54, 54, 54, 54, 54, 54, 54, 54, 54, 54, 54, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 55, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 56, 57, 57, 57, 57, 57, 57, 57, 57, 57, 57, 57, 57, 57, 57, 57, 57, 57, 57, 57, 57, 57, 57, 57, 57, 57, 57, 57, 57, 57, 57, 57, 57, 57, 57, 57, 57, 58, 58, 58, 58, 58, 58, 58, 58, 58, 58, 58, 58, 58, 58, 58, 58, 58, 58, 58, 58, 58, 58, 58, 58, 58, 58, 58, 58, 58, 58, 58, 58, 58, 58, 58, 58, 59, 59, 59, 59, 59, 59, 59, 59, 59, 59, 59, 59, 59, 59, 59, 59, 59, 59, 59, 59, 59, 59, 59, 59, 59, 59, 59, 59, 59, 59, 59, 59, 59, 59, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 60, 61, 61, 61, 61, 61, 61, 61, 61, 61, 61, 61, 61, 61, 61, 61, 61, 61, 61, 61, 61, 61, 61, 61, 61, 61, 61, 61, 61, 61, 61, 61, 61, 61, 62, 62, 62, 62, 62, 62, 62, 62, 62, 62, 62, 62, 62, 62, 62, 62, 62, 62, 62, 62, 62, 62, 62, 62, 62, 62, 62, 62, 62, 62, 62, 62, 62, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 63, 64, 64, 64, 64, 64, 64, 64, 64, 64, 64, 64, 64, 64, 64, 64, 64, 64, 64, 64, 64, 64, 64, 64, 64, 64, 64, 64, 64, 64, 64, 64, 64, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 65, 66, 66, 66, 66, 66, 66, 66, 66, 66, 66, 66, 66, 66, 66, 66, 66, 66, 66, 66, 66, 66, 66, 66, 66, 66, 66, 66, 66, 66, 66, 66, 67, 67, 67, 67, 67, 67, 67, 67, 67, 67, 67, 67, 67, 67, 67, 67, 67, 67, 67, 67, 67, 67, 67, 67, 67, 67, 67, 67, 67, 67, 67, 68, 68, 68, 68, 68, 68, 68, 68, 68, 68, 68, 68, 68, 68, 68, 68, 68, 68, 68, 68, 68, 68, 68, 68, 68, 68, 68, 68, 68, 68, 69, 69, 69, 69, 69, 69, 69, 69, 69, 69, 69, 69, 69, 69, 69, 69, 69, 69, 69, 69, 69, 69, 69, 69, 69, 69, 69, 69, 69, 69, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 70, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 71, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 72, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 73, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 74, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 75, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 76, 77, 77, 77, 77, 77, 77, 77, 77, 77, 77, 77, 77, 77, 77, 77, 77, 77, 77, 77, 77, 77, 77, 77, 77, 77, 77, 78, 78, 78, 78, 78, 78, 78, 78, 78, 78, 78, 78, 78, 78, 78, 78, 78, 78, 78, 78, 78, 78, 78, 78, 78, 78, 78, 79, 79, 79, 79, 79, 79, 79, 79, 79, 79, 79, 79, 79, 79, 79, 79, 79, 79, 79, 79, 79, 79, 79, 79, 79, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 80, 81, 81, 81, 81, 81, 81, 81, 81, 81, 81, 81, 81, 81, 81, 81, 81, 81, 81, 81, 81, 81, 81, 81, 81, 81, 82, 82, 82, 82, 82, 82, 82, 82, 82, 82, 82, 82, 82, 82, 82, 82, 82, 82, 82, 82, 82, 82, 82, 82, 82, 83, 83, 83, 83, 83, 83, 83, 83, 83, 83, 83, 83, 83, 83, 83, 83, 83, 83, 83, 83, 83, 83, 83, 83, 83, 84, 84, 84, 84, 84, 84, 84, 84, 84, 84, 84, 84, 84, 84, 84, 84, 84, 84, 84, 84, 84, 84, 84, 84, 84, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 85, 86, 86, 86, 86, 86, 86, 86, 86, 86, 86, 86, 86, 86, 86, 86, 86, 86, 86, 86, 86, 86, 86, 86, 86, 87, 87, 87, 87, 87, 87, 87, 87, 87, 87, 87, 87, 87, 87, 87, 87, 87, 87, 87, 87, 87, 87, 87, 88, 88, 88, 88, 88, 88, 88, 88, 88, 88, 88, 88, 88, 88, 88, 88, 88, 88, 88, 88, 88, 88, 88, 89, 89, 89, 89, 89, 89, 89, 89, 89, 89, 89, 89, 89, 89, 89, 89, 89, 89, 89, 89, 89, 89, 89, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 90, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 91, 92, 92, 92, 92, 92, 92, 92, 92, 92, 92, 92, 92, 92, 92, 92, 92, 92, 92, 92, 92, 92, 92, 93, 93, 93, 93, 93, 93, 93, 93, 93, 93, 93, 93, 93, 93, 93, 93, 93, 93, 93, 93, 93, 93, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 94, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 95, 96, 96, 96, 96, 96, 96, 96, 96, 96, 96, 96, 96, 96, 96, 96, 96, 96, 96, 96, 96, 96, 97, 97, 97, 97, 97, 97, 97, 97, 97, 97, 97, 97, 97, 97, 97, 97, 97, 97, 97, 97, 97, 98, 98, 98, 98, 98, 98, 98, 98, 98, 98, 98, 98, 98, 98, 98, 98, 98, 98, 98, 98, 98, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 99, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 100, 101, 101, 101, 101, 101, 101, 101, 101, 101, 101, 101, 101, 101, 101, 101, 101, 101, 101, 101, 101, 101, 102, 102, 102, 102, 102, 102, 102, 102, 102, 102, 102, 102, 102, 102, 102, 102, 102, 102, 102, 102, 103, 103, 103, 103, 103, 103, 103, 103, 103, 103, 103, 103, 103, 103, 103, 103, 103, 103, 103, 103, 104, 104, 104, 104, 104, 104, 104, 104, 104, 104, 104, 104, 104, 104, 104, 104, 104, 104, 104, 105, 105, 105, 105, 105, 105, 105, 105, 105, 105, 105, 105, 105, 105, 105, 105, 105, 105, 105, 105, 106, 106, 106, 106, 106, 106, 106, 106, 106, 106, 106, 106, 106, 106, 106, 106, 106, 106, 106, 107, 107, 107, 107, 107, 107, 107, 107, 107, 107, 107, 107, 107, 107, 107, 107, 107, 107, 107, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 108, 109, 109, 109, 109, 109, 109, 109, 109, 109, 109, 109, 109, 109, 109, 109, 109, 109, 109, 109, 110, 110, 110, 110, 110, 110, 110, 110, 110, 110, 110, 110, 110, 110, 110, 110, 110, 110, 110, 111, 111, 111, 111, 111, 111, 111, 111, 111, 111, 111, 111, 111, 111, 111, 111, 111, 111, 112, 112, 112, 112, 112, 112, 112, 112, 112, 112, 112, 112, 112, 112, 112, 112, 112, 112, 112, 113, 113, 113, 113, 113, 113, 113, 113, 113, 113, 113, 113, 113, 113, 113, 113, 113, 113, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 114, 115, 115, 115, 115, 115, 115, 115, 115, 115, 115, 115, 115, 115, 115, 115, 115, 115, 115, 116, 116, 116, 116, 116, 116, 116, 116, 116, 116, 116, 116, 116, 116, 116, 116, 116, 117, 117, 117, 117, 117, 117, 117, 117, 117, 117, 117, 117, 117, 117, 117, 117, 117, 117, 118, 118, 118, 118, 118, 118, 118, 118, 118, 118, 118, 118, 118, 118, 118, 118, 118, 119, 119, 119, 119, 119, 119, 119, 119, 119, 119, 119, 119, 119, 119, 119, 119, 119, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 120, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 121, 122, 122, 122, 122, 122, 122, 122, 122, 122, 122, 122, 122, 122, 122, 122, 122, 122, 123, 123, 123, 123, 123, 123, 123, 123, 123, 123, 123, 123, 123, 123, 123, 123, 123, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 124, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 125, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 126, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 127, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 128, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 129, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 130, 131, 131, 131, 131, 131, 131, 131, 131, 131, 131, 131, 131, 131, 131, 131, 131, 132, 132, 132, 132, 132, 132, 132, 132, 132, 132, 132, 132, 132, 132, 132, 133, 133, 133, 133, 133, 133, 133, 133, 133, 133, 133, 133, 133, 133, 133, 133, 134, 134, 134, 134, 134, 134, 134, 134, 134, 134, 134, 134, 134, 134, 134, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 135, 136, 136, 136, 136, 136, 136, 136, 136, 136, 136, 136, 136, 136, 136, 136, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 137, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 138, 139, 139, 139, 139, 139, 139, 139, 139, 139, 139, 139, 139, 139, 139, 139, 140, 140, 140, 140, 140, 140, 140, 140, 140, 140, 140, 140, 140, 140, 140, 141, 141, 141, 141, 141, 141, 141, 141, 141, 141, 141, 141, 141, 141, 142, 142, 142, 142, 142, 142, 142, 142, 142, 142, 142, 142, 142, 142, 142, 143, 143, 143, 143, 143, 143, 143, 143, 143, 143, 143, 143, 143, 143, 144, 144, 144, 144, 144, 144, 144, 144, 144, 144, 144, 144, 144, 144, 145, 145, 145, 145, 145, 145, 145, 145, 145, 145, 145, 145, 145, 145, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 146, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 147, 148, 148, 148, 148, 148, 148, 148, 148, 148, 148, 148, 148, 148, 148, 149, 149, 149, 149, 149, 149, 149, 149, 149, 149, 149, 149, 149, 149, 150, 150, 150, 150, 150, 150, 150, 150, 150, 150, 150, 150, 150, 150, 151, 151, 151, 151, 151, 151, 151, 151, 151, 151, 151, 151, 151, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 152, 153, 153, 153, 153, 153, 153, 153, 153, 153, 153, 153, 153, 153, 154, 154, 154, 154, 154, 154, 154, 154, 154, 154, 154, 154, 154, 154, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 155, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 156, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 157, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 158, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 159, 160, 160, 160, 160, 160, 160, 160, 160, 160, 160, 160, 160, 160, 161, 161, 161, 161, 161, 161, 161, 161, 161, 161, 161, 161, 161, 162, 162, 162, 162, 162, 162, 162, 162, 162, 162, 162, 162, 163, 163, 163, 163, 163, 163, 163, 163, 163, 163, 163, 163, 163, 164, 164, 164, 164, 164, 164, 164, 164, 164, 164, 164, 164, 165, 165, 165, 165, 165, 165, 165, 165, 165, 165, 165, 165, 165, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 166, 167, 167, 167, 167, 167, 167, 167, 167, 167, 167, 167, 167, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 168, 169, 169, 169, 169, 169, 169, 169, 169, 169, 169, 169, 169, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 170, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 171, 172, 172, 172, 172, 172, 172, 172, 172, 172, 172, 172, 172, 173, 173, 173, 173, 173, 173, 173, 173, 173, 173, 173, 173, 174, 174, 174, 174, 174, 174, 174, 174, 174, 174, 174, 174, 175, 175, 175, 175, 175, 175, 175, 175, 175, 175, 175, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 176, 177, 177, 177, 177, 177, 177, 177, 177, 177, 177, 177, 177, 178, 178, 178, 178, 178, 178, 178, 178, 178, 178, 178, 179, 179, 179, 179, 179, 179, 179, 179, 179, 179, 179, 179, 180, 180, 180, 180, 180, 180, 180, 180, 180, 180, 180, 181, 181, 181, 181, 181, 181, 181, 181, 181, 181, 181, 182, 182, 182, 182, 182, 182, 182, 182, 182, 182, 182, 182, 183, 183, 183, 183, 183, 183, 183, 183, 183, 183, 183, 184, 184, 184, 184, 184, 184, 184, 184, 184, 184, 184, 185, 185, 185, 185, 185, 185, 185, 185, 185, 185, 185, 186, 186, 186, 186, 186, 186, 186, 186, 186, 186, 186, 187, 187, 187, 187, 187, 187, 187, 187, 187, 187, 187, 188, 188, 188, 188, 188, 188, 188, 188, 188, 188, 188, 189, 189, 189, 189, 189, 189, 189, 189, 189, 189, 189, 190, 190, 190, 190, 190, 190, 190, 190, 190, 190, 190, 191, 191, 191, 191, 191, 191, 191, 191, 191, 191, 192, 192, 192, 192, 192, 192, 192, 192, 192, 192, 192, 193, 193, 193, 193, 193, 193, 193, 193, 193, 193, 193, 194, 194, 194, 194, 194, 194, 194, 194, 194, 194, 195, 195, 195, 195, 195, 195, 195, 195, 195, 195, 195, 196, 196, 196, 196, 196, 196, 196, 196, 196, 196, 197, 197, 197, 197, 197, 197, 197, 197, 197, 197, 197, 198, 198, 198, 198, 198, 198, 198, 198, 198, 198, 199, 199, 199, 199, 199, 199, 199, 199, 199, 199, 199, 200, 200, 200, 200, 200, 200, 200, 200, 200, 200, 201, 201, 201, 201, 201, 201, 201, 201, 201, 201, 202, 202, 202, 202, 202, 202, 202, 202, 202, 202, 203, 203, 203, 203, 203, 203, 203, 203, 203, 203, 204, 204, 204, 204, 204, 204, 204, 204, 204, 204, 205, 205, 205, 205, 205, 205, 205, 205, 205, 205, 206, 206, 206, 206, 206, 206, 206, 206, 206, 206, 207, 207, 207, 207, 207, 207, 207, 207, 207, 207, 208, 208, 208, 208, 208, 208, 208, 208, 208, 208, 209, 209, 209, 209, 209, 209, 209, 209, 209, 209, 210, 210, 210, 210, 210, 210, 210, 210, 210, 210, 211, 211, 211, 211, 211, 211, 211, 211, 211, 211, 212, 212, 212, 212, 212, 212, 212, 212, 212, 213, 213, 213, 213, 213, 213, 213, 213, 213, 213, 214, 214, 214, 214, 214, 214, 214, 214, 214, 215, 215, 215, 215, 215, 215, 215, 215, 215, 215, 216, 216, 216, 216, 216, 216, 216, 216, 216, 216, 217, 217, 217, 217, 217, 217, 217, 217, 217, 218, 218, 218, 218, 218, 218, 218, 218, 218, 219, 219, 219, 219, 219, 219, 219, 219, 219, 219, 220, 220, 220, 220, 220, 220, 220, 220, 220, 221, 221, 221, 221, 221, 221, 221, 221, 221, 222, 222, 222, 222, 222, 222, 222, 222, 222, 222, 223, 223, 223, 223, 223, 223, 223, 223, 223, 224, 224, 224, 224, 224, 224, 224, 224, 224, 225, 225, 225, 225, 225, 225, 225, 225, 225, 226, 226, 226, 226, 226, 226, 226, 226, 226, 227, 227, 227, 227, 227, 227, 227, 227, 227, 228, 228, 228, 228, 228, 228, 228, 228, 228, 229, 229, 229, 229, 229, 229, 229, 229, 229, 230, 230, 230, 230, 230, 230, 230, 230, 230, 231, 231, 231, 231, 231, 231, 231, 231, 231, 232, 232, 232, 232, 232, 232, 232, 232, 232, 233, 233, 233, 233, 233, 233, 233, 233, 233, 234, 234, 234, 234, 234, 234, 234, 234, 234, 235, 235, 235, 235, 235, 235, 235, 235, 236, 236, 236, 236, 236, 236, 236, 236, 236, 237, 237, 237, 237, 237, 237, 237, 237, 237, 238, 238, 238, 238, 238, 238, 238, 238, 239, 239, 239, 239, 239, 239, 239, 239, 239, 240, 240, 240, 240, 240, 240, 240, 240, 240, 241, 241, 241, 241, 241, 241, 241, 241, 242, 242, 242, 242, 242, 242, 242, 242, 242, 243, 243, 243, 243, 243, 243, 243, 243, 244, 244, 244, 244, 244, 244, 244, 244, 244, 245, 245, 245, 245, 245, 245, 245, 245, 246, 246, 246, 246, 246, 246, 246, 246, 247, 247, 247, 247, 247, 247, 247, 247, 247, 248, 248, 248, 248, 248, 248, 248, 248, 249, 249, 249, 249, 249, 249, 249, 249, 250, 250, 250, 250, 250, 250, 250, 250, 251, 251, 251, 251, 251, 251, 251, 251, 251, 252, 252, 252, 252, 252, 252, 252, 252, 253, 253, 253, 253, 253, 253, 253, 253, 254, 254, 254, 254, 254, 254, 254, 254, 255, 255, 255, 255, 255, 255, 255, 255, 256, 256, 256, 256, 256, 256, 256, 256, 257, 257, 257, 257, 257, 257, 257, 257, 258, 258, 258, 258, 258, 258, 258, 258, 259, 259, 259, 259, 259, 259, 259, 259, 260, 260, 260, 260, 260, 260, 260, 260, 261, 261, 261, 261, 261, 261, 261, 261, 262, 262, 262, 262, 262, 262, 262, 262, 263, 263, 263, 263, 263, 263, 263, 264, 264, 264, 264, 264, 264, 264, 264, 265, 265, 265, 265, 265, 265, 265, 265, 266, 266, 266, 266, 266, 266, 266, 266, 267, 267, 267, 267, 267, 267, 267, 268, 268, 268, 268, 268, 268, 268, 268, 269, 269, 269, 269, 269, 269, 269, 269, 270, 270, 270, 270, 270, 270, 270, 271, 271, 271, 271, 271, 271, 271, 271, 272, 272, 272, 272, 272, 272, 272, 273, 273, 273, 273, 273, 273, 273, 273, 274, 274, 274, 274, 274, 274, 274, 275, 275, 275, 275, 275, 275, 275, 275, 276, 276, 276, 276, 276, 276, 276, 277, 277, 277, 277, 277, 277, 277, 277, 278, 278, 278, 278, 278, 278, 278, 279, 279, 279, 279, 279, 279, 279, 279, 280, 280, 280, 280, 280, 280, 280, 281, 281, 281, 281, 281, 281, 281, 282, 282, 282, 282, 282, 282, 282, 282, 283, 283, 283, 283, 283, 283, 283, 284, 284, 284, 284, 284, 284, 284, 285, 285, 285, 285, 285, 285, 285, 286, 286, 286, 286, 286, 286, 286, 287, 287, 287, 287, 287, 287, 287, 287, 288, 288, 288, 288, 288, 288, 288, 289, 289, 289, 289, 289, 289, 289, 290, 290, 290, 290, 290, 290, 290, 291, 291, 291, 291, 291, 291, 291, 292, 292, 292, 292, 292, 292, 292, 293, 293, 293, 293, 293, 293, 293, 294, 294, 294, 294, 294, 294, 294, 295, 295, 295, 295, 295, 295, 295, 296, 296, 296, 296, 296, 296, 296, 297, 297, 297, 297, 297, 297, 297, 298, 298, 298, 298, 298, 298, 298, 299, 299, 299, 299, 299, 299, 299, 300, 300, 300, 300, 300, 300, 300, 301, 301, 301, 301, 301, 301, 302, 302, 302, 302, 302, 302, 302, 303, 303, 303, 303, 303, 303, 303, 304, 304, 304, 304, 304, 304, 304, 305, 305, 305, 305, 305, 305, 305, 306, 306, 306, 306, 306, 306, 307, 307, 307, 307, 307, 307, 307, 308, 308, 308, 308, 308, 308, 308, 309, 309, 309, 309, 309, 309, 310, 310, 310, 310, 310, 310, 310, 311, 311, 311, 311, 311, 311, 311, 312, 312, 312, 312, 312, 312, 313, 313, 313, 313, 313, 313, 313, 314, 314, 314, 314, 314, 314, 315, 315, 315, 315, 315, 315, 315, 316, 316, 316, 316, 316, 316, 317, 317, 317, 317, 317, 317, 317, 318, 318, 318, 318, 318, 318, 319, 319, 319, 319, 319, 319, 319, 320, 320, 320, 320, 320, 320, 321, 321, 321, 321, 321, 321, 321, 322, 322, 322, 322, 322, 322, 323, 323, 323, 323, 323, 323, 324, 324, 324, 324, 324, 324, 324, 325, 325, 325, 325, 325, 325, 326, 326, 326, 326, 326, 326, 327, 327, 327, 327, 327, 327, 327, 328, 328, 328, 328, 328, 328, 329, 329, 329, 329, 329, 329, 330, 330, 330, 330, 330, 330, 331, 331, 331, 331, 331, 331, 331, 332, 332, 332, 332, 332, 332, 333, 333, 333, 333, 333, 333, 334, 334, 334, 334, 334, 334, 335, 335, 335, 335, 335, 335, 336, 336, 336, 336, 336, 336, 337, 337, 337, 337, 337, 337, 337, 338, 338, 338, 338, 338, 338, 339, 339, 339, 339, 339, 339, 340, 340, 340, 340, 340, 340, 341, 341, 341, 341, 341, 341, 342, 342, 342, 342, 342, 342, 343, 343, 343, 343, 343, 343, 344, 344, 344, 344, 344, 344, 345, 345, 345, 345, 345, 345, 346, 346, 346, 346, 346, 346, 347, 347, 347, 347, 347, 347, 348, 348, 348, 348, 348, 348, 349, 349, 349, 349, 349, 349, 350, 350, 350, 350, 350, 351, 351, 351, 351, 351, 351, 352, 352, 352, 352, 352, 352, 353, 353, 353, 353, 353, 353, 354, 354, 354, 354, 354, 354, 355, 355, 355, 355, 355, 355, 356, 356, 356, 356, 356, 357, 357, 357, 357, 357, 357, 358, 358, 358, 358, 358, 358, 359, 359, 359, 359, 359, 359, 360, 360, 360, 360, 360, 361, 361, 361, 361, 361, 361, 362, 362, 362, 362, 362, 362, 363, 363, 363, 363, 363, 364, 364, 364, 364, 364, 364, 365, 365, 365, 365, 365, 365, 366, 366, 366, 366, 366, 367, 367, 367, 367, 367, 367, 368, 368, 368, 368, 368, 368, 369, 369, 369, 369, 369, 370, 370, 370, 370, 370, 370, 371, 371, 371, 371, 371, 372, 372, 372, 372, 372, 372, 373, 373, 373, 373, 373, 374, 374, 374, 374, 374, 374, 375, 375, 375, 375, 375, 376, 376, 376, 376, 376, 376, 377, 377, 377, 377, 377, 378, 378, 378, 378, 378, 378, 379, 379, 379, 379, 379, 380, 380, 380, 380, 380, 380, 381, 381, 381, 381, 381, 382, 382, 382, 382, 382, 383, 383, 383, 383, 383, 383, 384, 384, 384, 384, 384, 385, 385, 385, 385, 385, 386, 386, 386, 386, 386, 386, 387, 387, 387, 387, 387, 388, 388, 388, 388, 388, 389, 389, 389, 389, 389, 389, 390, 390, 390, 390, 390, 391, 391, 391, 391, 391, 392, 392, 392, 392, 392, 392, 393, 393, 393, 393, 393, 394, 394, 394, 394, 394, 395, 395, 395, 395, 395, 396, 396, 396, 396, 396, 397, 397, 397, 397, 397, 397, 398, 398, 398, 398, 398, 399, 399, 399, 399, 399, 400, 400, 400, 400, 400, 401, 401, 401, 401, 401, 402, 402, 402, 402, 402, 403, 403, 403, 403, 403, 404, 404, 404, 404, 404, 404, 405, 405, 405, 405, 405, 406, 406, 406, 406, 406, 407, 407, 407, 407, 407, 408, 408, 408, 408, 408, 409, 409, 409, 409, 409, 410, 410, 410, 410, 410, 411, 411, 411, 411, 411, 412, 412, 412, 412, 412, 413, 413, 413, 413, 413, 414, 414, 414, 414, 414, 415, 415, 415, 415, 415, 416, 416, 416, 416, 416, 417, 417, 417, 417, 417, 418, 418, 418, 418, 418, 419, 419, 419, 419, 419, 420, 420, 420, 420, 420, 421, 421, 421, 421, 422, 422, 422, 422, 422, 423, 423, 423, 423, 423, 424, 424, 424, 424, 424, 425, 425, 425, 425, 425, 426, 426, 426, 426, 426, 427, 427, 427, 427, 427, 428, 428, 428, 428, 429, 429, 429, 429, 429, 430, 430, 430, 430, 430, 431, 431, 431, 431, 431, 432, 432, 432, 432, 432, 433, 433, 433, 433, 434, 434, 434, 434, 434, 435, 435, 435, 435, 435, 436, 436, 436, 436, 437, 437, 437, 437, 437, 438, 438, 438, 438, 438, 439, 439, 439, 439, 439, 440, 440, 440, 440, 441, 441, 441, 441, 441, 442, 442, 442, 442, 442, 443, 443, 443, 443, 444, 444, 444, 444, 444, 445, 445, 445, 445, 445, 446, 446, 446, 446, 447, 447, 447, 447, 447, 448, 448, 448, 448, 449, 449, 449, 449, 449, 450, 450, 450, 450, 450, 451, 451, 451, 451, 452, 452, 452, 452, 452, 453, 453, 453, 453, 454, 454, 454, 454, 454, 455, 455, 455, 455, 456, 456, 456, 456, 456, 457, 457, 457, 457, 458, 458, 458, 458, 458, 459, 459, 459, 459, 460, 460, 460, 460, 460, 461, 461, 461, 461, 462, 462, 462, 462, 462, 463, 463, 463, 463, 464, 464, 464, 464, 464, 465, 465, 465, 465, 466, 466, 466, 466, 466, 467, 467, 467, 467, 468, 468, 468, 468, 469, 469, 469, 469, 469, 470, 470, 470, 470, 471, 471, 471, 471, 471, 472, 472, 472, 472, 473, 473, 473, 473, 474, 474, 474, 474, 474, 475, 475, 475, 475, 476, 476, 476, 476, 477, 477, 477, 477, 477, 478, 478, 478, 478, 479, 479, 479, 479, 480, 480, 480, 480, 480, 481, 481, 481, 481, 482, 482, 482, 482, 483, 483, 483, 483, 484, 484, 484, 484, 484, 485, 485, 485, 485, 486, 486, 486, 486, 487, 487, 487, 487, 488, 488, 488, 488, 488, 489, 489, 489, 489, 490, 490, 490, 490, 491, 491, 491, 491, 492, 492, 492, 492, 493, 493, 493, 493, 493, 494, 494, 494, 494, 495, 495, 495, 495, 496, 496, 496, 496, 497, 497, 497, 497, 498, 498, 498, 498, 499, 499, 499, 499, 499, 500, 500, 500, 500, 501, 501, 501, 501, 502, 502, 502, 502, 503, 503, 503, 503, 504, 504, 504, 504, 505, 505, 505, 505, 506, 506, 506, 506, 507, 507, 507, 507, 508, 508, 508, 508, 509, 509, 509, 509, 509, 510, 510, 510, 510, 511, 511, 511, 511, 512, 512, 512, 512, 513, 513, 513, 513, 514, 514, 514, 514, 515, 515, 515, 515, 516, 516, 516, 516, 517, 517, 517, 517, 518, 518, 518, 518, 519, 519, 519, 519, 520, 520, 520, 520, 521, 521, 521, 521, 522, 522, 522, 522, 523, 523, 523, 524, 524, 524, 524, 525, 525, 525, 525, 526, 526, 526, 526, 527, 527, 527, 527, 528, 528, 528, 528, 529, 529, 529, 529, 530, 530, 530, 530, 531, 531, 531, 531, 532, 532, 532, 532, 533, 533, 533, 533, 534, 534, 534, 535, 535, 535, 535, 536, 536, 536, 536, 537, 537, 537, 537, 538, 538, 538, 538, 539, 539, 539, 539, 540, 540, 540, 541, 541, 541, 541, 542, 542, 542, 542, 543, 543, 543, 543, 544, 544, 544, 544, 545, 545, 545, 546, 546, 546, 546, 547, 547, 547, 547, 548, 548, 548, 548, 549, 549, 549, 549, 550, 550, 550, 551, 551, 551, 551, 552, 552, 552, 552, 553, 553, 553, 553, 554, 554, 554, 555, 555, 555, 555, 556, 556, 556, 556, 557, 557, 557, 558, 558, 558, 558, 559, 559, 559, 559, 560, 560, 560, 561, 561, 561, 561, 562, 562, 562, 562, 563, 563, 563, 563, 564, 564, 564, 565, 565, 565, 565, 566, 566, 566, 567, 567, 567, 567, 568, 568, 568, 568, 569, 569, 569, 570, 570, 570, 570, 571, 571, 571, 571, 572, 572, 572, 573, 573, 573, 573, 574, 574, 574, 575, 575, 575, 575, 576, 576, 576, 576, 577, 577, 577, 578, 578, 578, 578, 579, 579, 579, 580, 580, 580, 580, 581, 581, 581, 582, 582, 582, 582, 583, 583, 583, 583, 584, 584, 584, 585, 585, 585, 585, 586, 586, 586, 587, 587, 587, 587, 588, 588, 588, 589, 589, 589, 589, 590, 590, 590, 591, 591, 591, 591, 592, 592, 592, 593, 593, 593, 593, 594, 594, 594, 595, 595, 595, 595, 596, 596, 596, 597, 597, 597, 597, 598, 598, 598, 599, 599, 599, 600, 600, 600, 600, 601, 601, 601, 602, 602, 602, 602, 603, 603, 603, 604, 604, 604, 604, 605, 605, 605, 606, 606, 606, 607, 607, 607, 607, 608, 608, 608, 609, 609, 609, 609, 610, 610, 610, 611, 611, 611, 612, 612, 612, 612, 613, 613, 613, 614, 614, 614, 614, 615, 615, 615, 616, 616, 616, 617, 617, 617, 617, 618, 618, 618, 619, 619, 619, 620, 620, 620, 620, 621, 621, 621, 622, 622, 622, 623, 623, 623, 623, 624, 624, 624, 625, 625, 625, 626, 626, 626, 626, 627, 627, 627, 628, 628, 628, 629, 629, 629, 630, 630, 630, 630, 631, 631, 631, 632, 632, 632, 633, 633, 633, 633, 634, 634, 634, 635, 635, 635, 636, 636, 636, 637, 637, 637, 637, 638, 638, 638, 639, 639, 639, 640, 640, 640, 641, 641, 641, 642, 642, 642, 642, 643, 643, 643, 644, 644, 644, 645, 645, 645, 646, 646, 646, 646, 647, 647, 647, 648, 648, 648, 649, 649, 649, 650, 650, 650, 651, 651, 651, 652, 652, 652, 652, 653, 653, 653, 654, 654, 654, 655, 655, 655, 656, 656, 656, 657, 657, 657, 658, 658, 658, 658, 659, 659, 659, 660, 660, 660, 661, 661, 661, 662, 662, 662, 663, 663, 663, 664, 664, 664, 665, 665, 665, 666, 666, 666, 666, 667, 667, 667, 668, 668, 668, 669, 669, 669, 670, 670, 670, 671, 671, 671, 672, 672, 672, 673, 673, 673, 674, 674, 674, 675, 675, 675, 676, 676, 676, 677, 677, 677, 678, 678, 678, 679, 679, 679, 679, 680, 680, 680, 681, 681, 681, 682, 682, 682, 683, 683, 683, 684, 684, 684, 685, 685, 685, 686, 686, 686, 687, 687, 687, 688, 688, 688, 689, 689, 689, 690, 690, 690, 691, 691, 691, 692, 692, 692, 693, 693, 693, 694, 694, 694, 695, 695, 695, 696, 696, 696, 697, 697, 697, 698, 698, 698, 699, 699, 699, 700, 700, 700, 701, 701, 702, 702, 702, 703, 703, 703, 704, 704, 704, 705, 705, 705, 706, 706, 706, 707, 707, 707, 708, 708, 708, 709, 709, 709, 710, 710, 710, 711, 711, 711, 712, 712, 712, 713, 713, 713, 714, 714, 714, 715, 715, 716, 716, 716, 717, 717, 717, 718, 718, 718, 719, 719, 719, 720, 720, 720, 721, 721, 721, 722, 722, 722, 723, 723, 724, 724, 724, 725, 725, 725, 726, 726, 726, 727, 727, 727, 728, 728, 728, 729, 729, 729, 730, 730, 731, 731, 731, 732, 732, 732, 733, 733, 733, 734, 734, 734, 735, 735, 736, 736, 736, 737, 737, 737, 738, 738, 738, 739, 739, 739, 740, 740, 740, 741, 741, 742, 742, 742, 743, 743, 743, 744, 744, 744, 745, 745, 746, 746, 746, 747, 747, 747, 748, 748, 748, 749, 749, 749, 750, 750, 751, 751, 751, 752, 752, 752, 753, 753, 753, 754, 754, 755, 755, 755, 756, 756, 756, 757, 757, 757, 758, 758, 759, 759, 759, 760, 760, 760, 761, 761, 762, 762, 762, 763, 763, 763, 764, 764, 764, 765, 765, 766, 766, 766, 767, 767, 767, 768, 768, 769, 769, 769, 770, 770, 770, 771, 771, 772, 772, 772, 773, 773, 773, 774, 774, 774, 775, 775, 776, 776, 776, 777, 777, 777, 778, 778, 779, 779, 779, 780, 780, 780, 781, 781, 782, 782, 782, 783, 783, 784, 784, 784, 785, 785, 785, 786, 786, 787, 787, 787, 788, 788, 788, 789, 789, 790, 790, 790, 791, 791, 791, 792, 792, 793, 793, 793, 794, 794, 795, 795, 795, 796, 796, 796, 797, 797, 798, 798, 798, 799, 799, 800, 800, 800, 801, 801, 801, 802, 802, 803, 803, 803, 804, 804, 805, 805, 805, 806, 806, 807, 807, 807, 808, 808, 808, 809, 809, 810, 810, 810, 811, 811, 812, 812, 812, 813, 813, 814, 814, 814, 815, 815, 816, 816, 816, 817, 817, 817, 818, 818, 819, 819, 819, 820, 820, 821, 821, 821, 822, 822, 823, 823, 823, 824, 824, 825, 825, 825, 826, 826, 827, 827, 827, 828, 828, 829, 829, 829, 830, 830, 831, 831, 831, 832, 832, 833, 833, 833, 834, 834, 835, 835, 835, 836, 836, 837, 837, 837, 838, 838, 839, 839, 839, 840, 840, 841, 841, 841, 842, 842, 843, 843, 843, 844, 844, 845, 845, 846, 846, 846, 847, 847, 848, 848, 848, 849, 849, 850, 850, 850, 851, 851, 852, 852, 852, 853, 853, 854, 854, 855, 855, 855, 856, 856, 857, 857, 857, 858, 858, 859, 859, 860, 860, 860, 861, 861, 862, 862, 862, 863, 863, 864, 864, 864, 865, 865, 866, 866, 867, 867, 867, 868, 868, 869, 869, 869, 870, 870, 871, 871, 872, 872, 872, 873, 873, 874, 874, 875, 875, 875, 876, 876, 877, 877, 877, 878, 878, 879, 879, 880, 880, 880, 881, 881, 882, 882, 883, 883, 883, 884, 884, 885, 885, 886, 886, 886, 887, 887, 888, 888, 889, 889, 889, 890, 890, 891, 891, 892, 892, 892, 893, 893, 894, 894, 895, 895, 895, 896, 896, 897, 897, 898, 898, 898, 899, 899, 900, 900, 901, 901, 901, 902, 902, 903, 903, 904, 904, 905, 905, 905, 906, 906, 907, 907, 908, 908, 908, 909, 909, 910, 910, 911, 911, 912, 912, 912, 913, 913, 914, 914, 915, 915, 915, 916, 916, 917, 917, 918, 918, 919, 919, 919, 920, 920, 921, 921, 922, 922, 923, 923, 923, 924, 924, 925, 925, 926, 926, 927, 927, 927, 928, 928, 929, 929, 930, 930, 931, 931, 931, 932, 932, 933, 933, 934, 934, 935, 935, 936, 936, 936, 937, 937, 938, 938, 939, 939, 940, 940, 940, 941, 941, 942, 942, 943, 943, 944, 944, 945, 945, 945, 946, 946, 947, 947, 948, 948, 949, 949, 950, 950, 951, 951, 951, 952, 952, 953, 953, 954, 954, 955, 955, 956, 956, 956, 957, 957, 958, 958, 959, 959, 960, 960, 961, 961, 962, 962, 962, 963, 963, 964, 964, 965, 965, 966, 966, 967, 967, 968, 968, 969, 969, 969, 970, 970, 971, 971, 972, 972, 973, 973, 974, 974, 975, 975, 976, 976, 976, 977, 977, 978, 978, 979, 979, 980, 980, 981, 981, 982, 982, 983, 983, 984, 984, 984, 985, 985, 986, 986, 987, 987, 988, 988, 989, 989, 990, 990, 991, 991, 992, 992, 993, 993, 994, 994, 994, 995, 995, 996, 996, 997, 997, 998, 998, 999, 999, 1000, 1000, 1001, 1001, 1002, 1002, 1003, 1003, 1004, 1004, 1005, 1005, 1006, 1006, 1006, 1007, 1007, 1008, 1008, 1009, 1009, 1010, 1010, 1011, 1011, 1012, 1012, 1013, 1013, 1014, 1014, 1015, 1015, 1016, 1016, 1017, 1017, 1018, 1018, 1019, 1019, 1020, 1020, 1021, 1021, 1022, 1022, 1023, 1023, 1024, 1024, 1025, 1025, 1026, 1026, 1027, 1027, 1028, 1028, 1029, 1029, 1029, 1030, 1030, 1031, 1031, 1032, 1032, 1033, 1033, 1034, 1034, 1035, 1035, 1036, 1036, 1037, 1037, 1038, 1038, 1039, 1039, 1040, 1040, 1041, 1041, 1042, 1042, 1043, 1043, 1044, 1044, 1045, 1045, 1046, 1046, 1047, 1047, 1048, 1048, 1049, 1049, 1050, 1050, 1051, 1051, 1052, 1053, 1053, 1054, 1054, 1055, 1055, 1056, 1056, 1057, 1057, 1058, 1058, 1059, 1059, 1060, 1060, 1061, 1061, 1062, 1062, 1063, 1063, 1064, 1064, 1065, 1065, 1066, 1066, 1067, 1067, 1068, 1068, 1069, 1069, 1070, 1070, 1071, 1071, 1072, 1072, 1073, 1073, 1074, 1074, 1075, 1076, 1076, 1077, 1077, 1078, 1078, 1079, 1079, 1080, 1080, 1081, 1081, 1082, 1082, 1083, 1083, 1084, 1084, 1085, 1085, 1086, 1086, 1087, 1087, 1088, 1088, 1089, 1090, 1090, 1091, 1091, 1092, 1092, 1093, 1093, 1094, 1094, 1095, 1095, 1096, 1096, 1097, 1097, 1098, 1098, 1099, 1100, 1100, 1101, 1101, 1102, 1102, 1103, 1103, 1104, 1104, 1105, 1105, 1106, 1106, 1107, 1107, 1108, 1109, 1109, 1110, 1110, 1111, 1111, 1112, 1112, 1113, 1113, 1114, 1114, 1115, 1115, 1116, 1117, 1117, 1118, 1118, 1119, 1119, 1120, 1120, 1121, 1121, 1122, 1122, 1123, 1124, 1124, 1125, 1125, 1126, 1126, 1127, 1127, 1128, 1128, 1129, 1129, 1130, 1131, 1131, 1132, 1132, 1133, 1133, 1134, 1134, 1135, 1135, 1136, 1137, 1137, 1138, 1138, 1139, 1139, 1140, 1140, 1141, 1141, 1142, 1143, 1143, 1144, 1144, 1145, 1145, 1146, 1146, 1147, 1148, 1148, 1149, 1149, 1150, 1150, 1151, 1151, 1152, 1152, 1153, 1154, 1154, 1155, 1155, 1156, 1156, 1157, 1157, 1158, 1159, 1159, 1160, 1160, 1161, 1161, 1162, 1162, 1163, 1164, 1164, 1165, 1165, 1166, 1166, 1167, 1167, 1168, 1169, 1169, 1170, 1170, 1171, 1171, 1172, 1173, 1173, 1174, 1174, 1175, 1175, 1176, 1176, 1177, 1178, 1178, 1179, 1179, 1180, 1180, 1181, 1182, 1182, 1183, 1183, 1184, 1184, 1185, 1186, 1186, 1187, 1187, 1188, 1188, 1189, 1190, 1190, 1191, 1191, 1192, 1192, 1193, 1194, 1194, 1195, 1195, 1196, 1196, 1197, 1198, 1198, 1199, 1199, 1200, 1200, 1201, 1202, 1202, 1203, 1203, 1204, 1204, 1205, 1206, 1206, 1207, 1207, 1208, 1208, 1209, 1210, 1210, 1211, 1211, 1212, 1213, 1213, 1214, 1214, 1215, 1215, 1216, 1217, 1217, 1218, 1218, 1219, 1220, 1220, 1221, 1221, 1222, 1222, 1223, 1224, 1224, 1225, 1225, 1226, 1227, 1227, 1228, 1228, 1229, 1230, 1230, 1231, 1231, 1232, 1232, 1233, 1234, 1234, 1235, 1235, 1236, 1237, 1237, 1238, 1238, 1239, 1240, 1240, 1241, 1241, 1242, 1243, 1243, 1244, 1244, 1245, 1246, 1246, 1247, 1247, 1248, 1249, 1249, 1250, 1250, 1251, 1252, 1252, 1253, 1253, 1254, 1255, 1255, 1256, 1256, 1257, 1258, 1258, 1259, 1259, 1260, 1261, 1261, 1262, 1262, 1263, 1264, 1264, 1265, 1265, 1266, 1267, 1267, 1268, 1268, 1269, 1270, 1270, 1271, 1271, 1272, 1273, 1273, 1274, 1274, 1275, 1276, 1276, 1277, 1278, 1278, 1279, 1279, 1280, 1281, 1281, 1282, 1282, 1283, 1284, 1284, 1285, 1286, 1286, 1287, 1287, 1288, 1289, 1289, 1290, 1290, 1291, 1292, 1292, 1293, 1294, 1294, 1295, 1295, 1296, 1297, 1297, 1298, 1299, 1299, 1300, 1300, 1301, 1302, 1302, 1303, 1303, 1304, 1305, 1305, 1306, 1307, 1307, 1308, 1308, 1309, 1310, 1310, 1311, 1312, 1312, 1313, 1314, 1314, 1315, 1315, 1316, 1317, 1317, 1318, 1319, 1319, 1320, 1320, 1321, 1322, 1322, 1323, 1324, 1324, 1325, 1326, 1326, 1327, 1327, 1328, 1329, 1329, 1330, 1331, 1331, 1332, 1333, 1333, 1334, 1334, 1335, 1336, 1336, 1337, 1338, 1338, 1339, 1340, 1340, 1341, 1341, 1342, 1343, 1343, 1344, 1345, 1345, 1346, 1347, 1347, 1348, 1349, 1349, 1350, 1350, 1351, 1352, 1352, 1353, 1354, 1354, 1355, 1356, 1356, 1357, 1358, 1358, 1359, 1360, 1360, 1361, 1361, 1362, 1363, 1363, 1364, 1365, 1365, 1366, 1367, 1367, 1368, 1369, 1369, 1370, 1371, 1371, 1372, 1373, 1373, 1374, 1375, 1375, 1376, 1377, 1377, 1378, 1379, 1379, 1380, 1380, 1381, 1382, 1382, 1383, 1384, 1384, 1385, 1386, 1386, 1387, 1388, 1388, 1389, 1390, 1390, 1391, 1392, 1392, 1393, 1394, 1394, 1395, 1396, 1396, 1397, 1398, 1398, 1399, 1400, 1400, 1401, 1402, 1402, 1403, 1404, 1404, 1405, 1406, 1406, 1407, 1408, 1408, 1409, 1410, 1411, 1411, 1412, 1413, 1413, 1414, 1415, 1415, 1416, 1417, 1417, 1418, 1419, 1419, 1420, 1421, 1421, 1422, 1423, 1423, 1424, 1425, 1425, 1426, 1427, 1427, 1428, 1429, 1429, 1430, 1431, 1432, 1432, 1433, 1434, 1434, 1435, 1436, 1436, 1437, 1438, 1438, 1439, 1440, 1440, 1441, 1442, 1443, 1443, 1444, 1445, 1445, 1446, 1447, 1447, 1448, 1449, 1449, 1450, 1451, 1452, 1452, 1453, 1454, 1454, 1455, 1456, 1456, 1457, 1458, 1458, 1459, 1460, 1461, 1461, 1462, 1463, 1463, 1464, 1465, 1465, 1466, 1467, 1468, 1468, 1469, 1470, 1470, 1471, 1472, 1472, 1473, 1474, 1475, 1475, 1476, 1477, 1477, 1478, 1479, 1479, 1480, 1481, 1482, 1482, 1483, 1484, 1484, 1485, 1486, 1487, 1487, 1488, 1489, 1489, 1490, 1491, 1492, 1492, 1493, 1494, 1494, 1495, 1496, 1497, 1497, 1498, 1499, 1499, 1500, 1501, 1502, 1502, 1503, 1504, 1504, 1505, 1506, 1507, 1507, 1508, 1509, 1509, 1510, 1511, 1512, 1512, 1513, 1514, 1514, 1515, 1516, 1517, 1517, 1518, 1519, 1520, 1520, 1521, 1522, 1522, 1523, 1524, 1525, 1525, 1526, 1527, 1528, 1528, 1529, 1530, 1530, 1531, 1532, 1533, 1533, 1534, 1535, 1536, 1536, 1537, 1538, 1539, 1539, 1540, 1541, 1541, 1542, 1543, 1544, 1544, 1545, 1546, 1547, 1547, 1548, 1549, 1550, 1550, 1551, 1552, 1553, 1553, 1554, 1555, 1555, 1556, 1557, 1558, 1558, 1559, 1560, 1561, 1561, 1562, 1563, 1564, 1564, 1565, 1566, 1567, 1567, 1568, 1569, 1570, 1570, 1571, 1572, 1573, 1573, 1574, 1575, 1576, 1576, 1577, 1578, 1579, 1579, 1580, 1581, 1582, 1582, 1583, 1584, 1585, 1585, 1586, 1587, 1588, 1588, 1589, 1590, 1591, 1591, 1592, 1593, 1594, 1595, 1595, 1596, 1597, 1598, 1598, 1599, 1600, 1601, 1601, 1602, 1603, 1604, 1604, 1605, 1606, 1607, 1607, 1608, 1609, 1610, 1611, 1611, 1612, 1613, 1614, 1614, 1615, 1616, 1617, 1617, 1618, 1619, 1620, 1621, 1621, 1622, 1623, 1624, 1624, 1625, 1626, 1627, 1627, 1628, 1629, 1630, 1631, 1631, 1632, 1633, 1634, 1634, 1635, 1636, 1637, 1638, 1638, 1639, 1640, 1641, 1642, 1642, 1643, 1644, 1645, 1645, 1646, 1647, 1648, 1649, 1649, 1650, 1651, 1652, 1652, 1653, 1654, 1655, 1656, 1656, 1657, 1658, 1659, 1660, 1660, 1661, 1662, 1663, 1664, 1664, 1665, 1666, 1667, 1667, 1668, 1669, 1670, 1671, 1671, 1672, 1673, 1674, 1675, 1675, 1676, 1677, 1678, 1679, 1679, 1680, 1681, 1682, 1683, 1683, 1684, 1685, 1686, 1687, 1687, 1688, 1689, 1690, 1691, 1691, 1692, 1693, 1694, 1695, 1695, 1696, 1697, 1698, 1699, 1700, 1700, 1701, 1702, 1703, 1704, 1704, 1705, 1706, 1707, 1708, 1708, 1709, 1710, 1711, 1712, 1713, 1713, 1714, 1715, 1716, 1717, 1717, 1718, 1719, 1720, 1721, 1721, 1722, 1723, 1724, 1725, 1726, 1726, 1727, 1728, 1729, 1730, 1731, 1731, 1732, 1733, 1734, 1735, 1735, 1736, 1737, 1738, 1739, 1740, 1740, 1741, 1742, 1743, 1744, 1745, 1745, 1746, 1747, 1748, 1749, 1750, 1750, 1751, 1752, 1753, 1754, 1755, 1755, 1756, 1757, 1758, 1759, 1760, 1760, 1761, 1762, 1763, 1764, 1765, 1765, 1766, 1767, 1768, 1769, 1770, 1770, 1771, 1772, 1773, 1774, 1775, 1775, 1776, 1777, 1778, 1779, 1780, 1781, 1781, 1782, 1783, 1784, 1785, 1786, 1786, 1787, 1788, 1789, 1790, 1791, 1792, 1792, 1793, 1794, 1795, 1796, 1797, 1798, 1798, 1799, 1800, 1801, 1802, 1803, 1804, 1804, 1805, 1806, 1807, 1808, 1809, 1810, 1810, 1811, 1812, 1813, 1814, 1815, 1816, 1816, 1817, 1818, 1819, 1820, 1821, 1822, 1822, 1823, 1824, 1825, 1826, 1827, 1828, 1829, 1829, 1830, 1831, 1832, 1833, 1834, 1835, 1836, 1836, 1837, 1838, 1839, 1840, 1841, 1842, 1842, 1843, 1844, 1845, 1846, 1847, 1848, 1849, 1849, 1850, 1851, 1852, 1853, 1854, 1855, 1856, 1857, 1857, 1858, 1859, 1860, 1861, 1862, 1863, 1864, 1864, 1865, 1866, 1867, 1868, 1869, 1870, 1871, 1872, 1872, 1873, 1874, 1875, 1876, 1877, 1878, 1879, 1880, 1880, 1881, 1882, 1883, 1884, 1885, 1886, 1887, 1888, 1888, 1889, 1890, 1891, 1892, 1893, 1894, 1895, 1896, 1897, 1897, 1898, 1899, 1900, 1901, 1902, 1903, 1904, 1905, 1906, 1906, 1907, 1908, 1909, 1910, 1911, 1912, 1913, 1914, 1915, 1916, 1916, 1917, 1918, 1919, 1920, 1921, 1922, 1923, 1924, 1925, 1926, 1926, 1927, 1928, 1929, 1930, 1931, 1932, 1933, 1934, 1935, 1936, 1937, 1937, 1938, 1939, 1940, 1941, 1942, 1943, 1944, 1945, 1946, 1947, 1948, 1949, 1949, 1950, 1951, 1952, 1953, 1954, 1955, 1956, 1957, 1958, 1959, 1960, 1961, 1961, 1962, 1963, 1964, 1965, 1966, 1967, 1968, 1969, 1970, 1971, 1972, 1973, 1974, 1975, 1975, 1976, 1977, 1978, 1979, 1980, 1981, 1982, 1983, 1984, 1985, 1986, 1987, 1988, 1989, 1990, 1990, 1991, 1992, 1993, 1994, 1995, 1996, 1997, 1998, 1999, 2000, 2001, 2002, 2003, 2004, 2005, 2006, 2007, 2008, 2008, 2009, 2010, 2011, 2012, 2013, 2014, 2015, 2016, 2017, 2018, 2019, 2020, 2021, 2022, 2023, 2024, 2025, 2026, 2027, 2028, 2029, 2029, 2030, 2031, 2032, 2033, 2034, 2035, 2036, 2037, 2038, 2039, 2040, 2041, 2042, 2043, 2044, 2045, 2046, 2047, 2048, 2049, 2050, 2051, 2052, 2053, 2054, 2055, 2056, 2057, 2058, 2058, 2059, 2060, 2061, 2062, 2063, 2064, 2065, 2066, 2067, 2068, 2069, 2070, 2071, 2072, 2073, 2074, 2075, 2076, 2077, 2078, 2079, 2080, 2081, 2082, 2083, 2084, 2085, 2086, 2087, 2088, 2089, 2090, 2091, 2092, 2093, 2094, 2095, 2096, 2097, 2098, 2099, 2100, 2101, 2102, 2103, 2104, 2105, 2106, 2107, 2108, 2109, 2110, 2111, 2112, 2113, 2114, 2115, 2116, 2117, 2118, 2119, 2120, 2121, 2122, 2123, 2124, 2125, 2126, 2127, 2128, 2129, 2130, 2131, 2132, 2133, 2134, 2135, 2136, 2137, 2138, 2139, 2140, 2141, 2142, 2143, 2144, 2145, 2146, 2147, 2148, 2149, 2150, 2151, 2152, 2153, 2154, 2155, 2156, 2157, 2158, 2159, 2160, 2161, 2162, 2163, 2164, 2165, 2166, 2167, 2168, 2169, 2170, 2171, 2172, 2173, 2174, 2176, 2177, 2178, 2179, 2180, 2181, 2182, 2183, 2184, 2185, 2186, 2187, 2188, 2189, 2190, 2191, 2192, 2193, 2194, 2195, 2196, 2197, 2198, 2199, 2200, 2201, 2202, 2203, 2204, 2205, 2207, 2208, 2209, 2210, 2211, 2212, 2213, 2214, 2215, 2216, 2217, 2218, 2219, 2220, 2221, 2222, 2223, 2224, 2225, 2226, 2227, 2228, 2230, 2231, 2232, 2233, 2234, 2235, 2236, 2237, 2238, 2239, 2240, 2241, 2242, 2243, 2244, 2245, 2246, 2247, 2249, 2250, 2251, 2252, 2253, 2254, 2255, 2256, 2257, 2258, 2259, 2260, 2261, 2262, 2263, 2265, 2266, 2267, 2268, 2269, 2270, 2271, 2272, 2273, 2274, 2275, 2276, 2277, 2278, 2279, 2281, 2282, 2283, 2284, 2285, 2286, 2287, 2288, 2289, 2290, 2291, 2292, 2294, 2295, 2296, 2297, 2298, 2299, 2300, 2301, 2302, 2303, 2304, 2305, 2307, 2308, 2309, 2310, 2311, 2312, 2313, 2314, 2315, 2316, 2317, 2318, 2320, 2321, 2322, 2323, 2324, 2325, 2326, 2327, 2328, 2329, 2331, 2332, 2333, 2334, 2335, 2336, 2337, 2338, 2339, 2340, 2342, 2343, 2344, 2345, 2346, 2347, 2348, 2349, 2350, 2351, 2353, 2354, 2355, 2356, 2357, 2358, 2359, 2360, 2361, 2363, 2364, 2365, 2366, 2367, 2368, 2369, 2370, 2371, 2373, 2374, 2375, 2376, 2377, 2378, 2379, 2380, 2382, 2383, 2384, 2385, 2386, 2387, 2388, 2389, 2391, 2392, 2393, 2394, 2395, 2396, 2397, 2398, 2400, 2401, 2402, 2403, 2404, 2405, 2406, 2407, 2409, 2410, 2411, 2412, 2413, 2414, 2415, 2417, 2418, 2419, 2420, 2421, 2422, 2423, 2425, 2426, 2427, 2428, 2429, 2430, 2431, 2432, 2434, 2435, 2436, 2437, 2438, 2439, 2441, 2442, 2443, 2444, 2445, 2446, 2447, 2449, 2450, 2451, 2452, 2453, 2454, 2455, 2457, 2458, 2459, 2460, 2461, 2462, 2464, 2465, 2466, 2467, 2468, 2469, 2471, 2472, 2473, 2474, 2475, 2476, 2477, 2479, 2480, 2481, 2482, 2483, 2484, 2486, 2487, 2488, 2489, 2490, 2491, 2493, 2494, 2495, 2496, 2497, 2499, 2500, 2501, 2502, 2503, 2504, 2506, 2507, 2508, 2509, 2510, 2511, 2513, 2514, 2515, 2516, 2517, 2519, 2520, 2521, 2522, 2523, 2524, 2526, 2527, 2528, 2529, 2530, 2532, 2533, 2534, 2535, 2536, 2538, 2539, 2540, 2541, 2542, 2544, 2545, 2546, 2547, 2548, 2549, 2551, 2552, 2553, 2554, 2555, 2557, 2558, 2559, 2560, 2561, 2563, 2564, 2565, 2566, 2567, 2569, 2570, 2571, 2572, 2574, 2575, 2576, 2577, 2578, 2580, 2581, 2582, 2583, 2584, 2586, 2587, 2588, 2589, 2590, 2592, 2593, 2594, 2595, 2597, 2598, 2599, 2600, 2601, 2603, 2604, 2605, 2606, 2608, 2609, 2610, 2611, 2612, 2614, 2615, 2616, 2617, 2619, 2620, 2621, 2622, 2623, 2625, 2626, 2627, 2628, 2630, 2631, 2632, 2633, 2635, 2636, 2637, 2638, 2640, 2641, 2642, 2643, 2644, 2646, 2647, 2648, 2649, 2651, 2652, 2653, 2654, 2656, 2657, 2658, 2659, 2661, 2662, 2663, 2664, 2666, 2667, 2668, 2669, 2671, 2672, 2673, 2674, 2676, 2677, 2678, 2679, 2681, 2682, 2683, 2684, 2686, 2687, 2688, 2689, 2691, 2692, 2693, 2694, 2696, 2697, 2698, 2700, 2701, 2702, 2703, 2705, 2706, 2707, 2708, 2710, 2711, 2712, 2713, 2715, 2716, 2717, 2719, 2720, 2721, 2722, 2724, 2725, 2726, 2727, 2729, 2730, 2731, 2733, 2734, 2735, 2736, 2738, 2739, 2740, 2742, 2743, 2744, 2745, 2747, 2748, 2749, 2751, 2752, 2753, 2754, 2756, 2757, 2758, 2760, 2761, 2762, 2763, 2765, 2766, 2767, 2769, 2770, 2771, 2772, 2774, 2775, 2776, 2778, 2779, 2780, 2782, 2783, 2784, 2785, 2787, 2788, 2789, 2791, 2792, 2793, 2795, 2796, 2797, 2799, 2800, 2801, 2802, 2804, 2805, 2806, 2808, 2809, 2810, 2812, 2813, 2814, 2816, 2817, 2818, 2820, 2821, 2822, 2823, 2825, 2826, 2827, 2829, 2830, 2831, 2833, 2834, 2835, 2837, 2838, 2839, 2841, 2842, 2843, 2845, 2846, 2847, 2849, 2850, 2851, 2853, 2854, 2855, 2857, 2858, 2859, 2861, 2862, 2863, 2865, 2866, 2867, 2869, 2870, 2871, 2873, 2874, 2875, 2877, 2878, 2879, 2881, 2882, 2883, 2885, 2886, 2888, 2889, 2890, 2892, 2893, 2894, 2896, 2897, 2898, 2900, 2901, 2902, 2904, 2905, 2906, 2908, 2909, 2910, 2912, 2913, 2915, 2916, 2917, 2919, 2920, 2921, 2923, 2924, 2925, 2927, 2928, 2930, 2931, 2932, 2934, 2935, 2936, 2938, 2939, 2941, 2942, 2943, 2945, 2946, 2947, 2949, 2950, 2952, 2953, 2954, 2956, 2957, 2958, 2960, 2961, 2963, 2964, 2965, 2967, 2968, 2969, 2971, 2972, 2974, 2975, 2976, 2978, 2979, 2981, 2982, 2983, 2985, 2986, 2988, 2989, 2990, 2992, 2993, 2994, 2996, 2997, 2999, 3000, 3001, 3003, 3004, 3006, 3007, 3008, 3010, 3011, 3013, 3014, 3015, 3017, 3018, 3020, 3021, 3023, 3024, 3025, 3027, 3028, 3030, 3031, 3032, 3034, 3035, 3037, 3038, 3039, 3041, 3042, 3044, 3045, 3047, 3048, 3049, 3051, 3052, 3054, 3055, 3056, 3058, 3059, 3061, 3062, 3064, 3065, 3066, 3068, 3069, 3071, 3072, 3074, 3075, 3076, 3078, 3079, 3081, 3082, 3084, 3085, 3086, 3088, 3089, 3091, 3092, 3094, 3095, 3097, 3098, 3099, 3101, 3102, 3104, 3105, 3107, 3108, 3110, 3111, 3112, 3114, 3115, 3117, 3118, 3120, 3121, 3123, 3124, 3125, 3127, 3128, 3130, 3131, 3133, 3134, 3136, 3137, 3139, 3140, 3142, 3143, 3144, 3146, 3147, 3149, 3150, 3152, 3153, 3155, 3156, 3158, 3159, 3161, 3162, 3164, 3165, 3166, 3168, 3169, 3171, 3172, 3174, 3175, 3177, 3178, 3180, 3181, 3183, 3184, 3186, 3187, 3189, 3190, 3192, 3193, 3195, 3196, 3197, 3199, 3200, 3202, 3203, 3205, 3206, 3208, 3209, 3211, 3212, 3214, 3215, 3217, 3218, 3220, 3221, 3223, 3224, 3226, 3227, 3229, 3230, 3232, 3233, 3235, 3236, 3238, 3239, 3241, 3242, 3244, 3245, 3247, 3248, 3250, 3251, 3253, 3254, 3256, 3257, 3259, 3260, 3262, 3263, 3265, 3266, 3268, 3270, 3271, 3273, 3274, 3276, 3277, 3279, 3280, 3282, 3283, 3285, 3286, 3288, 3289, 3291, 3292, 3294, 3295, 3297, 3298, 3300, 3302, 3303, 3305, 3306, 3308, 3309, 3311, 3312, 3314, 3315, 3317, 3318, 3320, 3321, 3323, 3325, 3326, 3328, 3329, 3331, 3332, 3334, 3335, 3337, 3338, 3340, 3342, 3343, 3345, 3346, 3348, 3349, 3351, 3352, 3354, 3356, 3357, 3359, 3360, 3362, 3363, 3365, 3366, 3368, 3370, 3371, 3373, 3374, 3376, 3377, 3379, 3380, 3382, 3384, 3385, 3387, 3388, 3390, 3391, 3393, 3395, 3396, 3398, 3399, 3401, 3402, 3404, 3406, 3407, 3409, 3410, 3412, 3414, 3415, 3417, 3418, 3420, 3421, 3423, 3425, 3426, 3428, 3429, 3431, 3433, 3434, 3436, 3437, 3439, 3440, 3442, 3444, 3445, 3447, 3448, 3450, 3452, 3453, 3455, 3456, 3458, 3460, 3461, 3463, 3464, 3466, 3468, 3469, 3471, 3472, 3474, 3476, 3477, 3479, 3480, 3482, 3484, 3485, 3487, 3489, 3490, 3492, 3493, 3495, 3497, 3498, 3500, 3501, 3503, 3505, 3506, 3508, 3510, 3511, 3513, 3514, 3516, 3518, 3519, 3521, 3523, 3524, 3526, 3527, 3529, 3531, 3532, 3534, 3536, 3537, 3539, 3541, 3542, 3544, 3545, 3547, 3549, 3550, 3552, 3554, 3555, 3557, 3559, 3560, 3562, 3563, 3565, 3567, 3568, 3570, 3572, 3573, 3575, 3577, 3578, 3580, 3582, 3583, 3585, 3587, 3588, 3590, 3592, 3593, 3595, 3597, 3598, 3600, 3602, 3603, 3605, 3606, 3608, 3610, 3611, 3613, 3615, 3616, 3618, 3620, 3621, 3623, 3625, 3627, 3628, 3630, 3632, 3633, 3635, 3637, 3638, 3640, 3642, 3643, 3645, 3647, 3648, 3650, 3652, 3653, 3655, 3657, 3658, 3660, 3662, 3663, 3665, 3667, 3669, 3670, 3672, 3674, 3675, 3677, 3679, 3680, 3682, 3684, 3686, 3687, 3689, 3691, 3692, 3694, 3696, 3697, 3699, 3701, 3703, 3704, 3706, 3708, 3709, 3711, 3713, 3714, 3716, 3718, 3720, 3721, 3723, 3725, 3726, 3728, 3730, 3732, 3733, 3735, 3737, 3739, 3740, 3742, 3744, 3745, 3747, 3749, 3751, 3752, 3754, 3756, 3757, 3759, 3761, 3763, 3764, 3766, 3768, 3770, 3771, 3773, 3775, 3777, 3778, 3780, 3782, 3784, 3785, 3787, 3789, 3790, 3792, 3794, 3796, 3797, 3799, 3801, 3803, 3804, 3806, 3808, 3810, 3811, 3813, 3815, 3817, 3818, 3820, 3822, 3824, 3826, 3827, 3829, 3831, 3833, 3834, 3836, 3838, 3840, 3841, 3843, 3845, 3847, 3848, 3850, 3852, 3854, 3856, 3857, 3859, 3861, 3863, 3864, 3866, 3868, 3870, 3871, 3873, 3875, 3877, 3879, 3880, 3882, 3884, 3886, 3888, 3889, 3891, 3893, 3895, 3896, 3898, 3900, 3902, 3904, 3905, 3907, 3909, 3911, 3913, 3914, 3916, 3918, 3920, 3922, 3923, 3925, 3927, 3929, 3931, 3932, 3934, 3936, 3938, 3940, 3941, 3943, 3945, 3947, 3949, 3951, 3952, 3954, 3956, 3958, 3960, 3961, 3963, 3965, 3967, 3969, 3970, 3972, 3974, 3976, 3978, 3980, 3981, 3983, 3985, 3987, 3989, 3991, 3992, 3994, 3996, 3998, 4000, 4002, 4003, 4005, 4007, 4009, 4011, 4013, 4014, 4016, 4018, 4020, 4022, 4024, 4025, 4027, 4029, 4031, 4033, 4035, 4037, 4038, 4040, 4042, 4044, 4046, 4048, 4050, 4051, 4053, 4055, 4057, 4059, 4061, 4063, 4064, 4066, 4068, 4070, 4072, 4074, 4076, 4077, 4079, 4081, 4083, 4085, 4087, 4089, 4091, 4092, 4094, 4096, 4098, 4100, 4102, 4104, 4106, 4107, 4109, 4111, 4113, 4115, 4117, 4119, 4121, 4122, 4124, 4126, 4128, 4130, 4132, 4134, 4136, 4138, 4140, 4141, 4143, 4145, 4147, 4149, 4151, 4153, 4155, 4157, 4158, 4160, 4162, 4164, 4166, 4168, 4170, 4172, 4174, 4176, 4178, 4179, 4181, 4183, 4185, 4187, 4189, 4191, 4193, 4195, 4197, 4199, 4201, 4202, 4204, 4206, 4208, 4210, 4212, 4214, 4216, 4218, 4220, 4222, 4224, 4226, 4227, 4229, 4231, 4233, 4235, 4237, 4239, 4241, 4243, 4245, 4247, 4249, 4251, 4253, 4255, 4257, 4258, 4260, 4262, 4264, 4266, 4268, 4270, 4272, 4274, 4276, 4278, 4280, 4282, 4284, 4286, 4288, 4290, 4292, 4294, 4296, 4298, 4299, 4301, 4303, 4305, 4307, 4309, 4311, 4313, 4315, 4317, 4319, 4321, 4323, 4325, 4327, 4329, 4331, 4333, 4335, 4337, 4339, 4341, 4343, 4345, 4347, 4349, 4351, 4353, 4355, 4357, 4359, 4361, 4363, 4365, 4367, 4369, 4371, 4373, 4375, 4377, 4379, 4381, 4383, 4385, 4387, 4389, 4391, 4393, 4395, 4397, 4399, 4401, 4403, 4405, 4407, 4409, 4411, 4413, 4415, 4417, 4419, 4421, 4423, 4425, 4427, 4429, 4431, 4433, 4435, 4437, 4439, 4441, 4443, 4445, 4447, 4449, 4451, 4453, 4455, 4457, 4459, 4461, 4463, 4465, 4467, 4469, 4471, 4473, 4475, 4477, 4479, 4481, 4484, 4486, 4488, 4490, 4492, 4494, 4496, 4498, 4500, 4502, 4504, 4506, 4508, 4510, 4512, 4514, 4516, 4518, 4520, 4522, 4524, 4527, 4529, 4531, 4533, 4535, 4537, 4539, 4541, 4543, 4545, 4547, 4549, 4551, 4553, 4555, 4557, 4560, 4562, 4564, 4566, 4568, 4570, 4572, 4574, 4576, 4578, 4580, 4582, 4584, 4587, 4589, 4591, 4593, 4595, 4597, 4599, 4601, 4603, 4605, 4607, 4610, 4612, 4614, 4616, 4618, 4620, 4622, 4624, 4626, 4628, 4630, 4633, 4635, 4637, 4639, 4641, 4643, 4645, 4647, 4649, 4652, 4654, 4656, 4658, 4660, 4662, 4664, 4666, 4668, 4671, 4673, 4675, 4677, 4679, 4681, 4683, 4685, 4688, 4690, 4692, 4694, 4696, 4698, 4700, 4702, 4705, 4707, 4709, 4711, 4713, 4715, 4717, 4720, 4722, 4724, 4726, 4728, 4730, 4732, 4735, 4737, 4739, 4741, 4743, 4745, 4747, 4750, 4752, 4754, 4756, 4758, 4760, 4762, 4765, 4767, 4769, 4771, 4773, 4775, 4778, 4780, 4782, 4784, 4786, 4788, 4791, 4793, 4795, 4797, 4799, 4801, 4804, 4806, 4808, 4810, 4812, 4814, 4817, 4819, 4821, 4823, 4825, 4828, 4830, 4832, 4834, 4836, 4839, 4841, 4843, 4845, 4847, 4849, 4852, 4854, 4856, 4858, 4860, 4863, 4865, 4867, 4869, 4871, 4874, 4876, 4878, 4880, 4882, 4885, 4887, 4889, 4891, 4893, 4896, 4898, 4900, 4902, 4905, 4907, 4909, 4911, 4913, 4916, 4918, 4920, 4922, 4925, 4927, 4929, 4931, 4933, 4936, 4938, 4940, 4942, 4945, 4947, 4949, 4951, 4954, 4956, 4958, 4960, 4962, 4965, 4967, 4969, 4971, 4974, 4976, 4978, 4980, 4983, 4985, 4987, 4989, 4992, 4994, 4996, 4998, 5001, 5003, 5005, 5007, 5010, 5012, 5014, 5016, 5019, 5021, 5023, 5026, 5028, 5030, 5032, 5035, 5037, 5039, 5041, 5044, 5046, 5048, 5051, 5053, 5055, 5057, 5060, 5062, 5064, 5066, 5069, 5071, 5073, 5076, 5078, 5080, 5082, 5085, 5087, 5089, 5092, 5094, 5096, 5099, 5101, 5103, 5105, 5108, 5110, 5112, 5115, 5117, 5119, 5122, 5124, 5126, 5128, 5131, 5133, 5135, 5138, 5140, 5142, 5145, 5147, 5149, 5152, 5154, 5156, 5159, 5161, 5163, 5166, 5168, 5170, 5172, 5175, 5177, 5179, 5182, 5184, 5186, 5189, 5191, 5193, 5196, 5198, 5200, 5203, 5205, 5207, 5210, 5212, 5215, 5217, 5219, 5222, 5224, 5226, 5229, 5231, 5233, 5236, 5238, 5240, 5243, 5245, 5247, 5250, 5252, 5254, 5257, 5259, 5262, 5264, 5266, 5269, 5271, 5273, 5276, 5278, 5281, 5283, 5285, 5288, 5290, 5292, 5295, 5297, 5300, 5302, 5304, 5307, 5309, 5311, 5314, 5316, 5319, 5321, 5323, 5326, 5328, 5331, 5333, 5335, 5338, 5340, 5342, 5345, 5347, 5350, 5352, 5354, 5357, 5359, 5362, 5364, 5366, 5369, 5371, 5374, 5376, 5379, 5381, 5383, 5386, 5388, 5391, 5393, 5395, 5398, 5400, 5403, 5405, 5408, 5410, 5412, 5415, 5417, 5420, 5422, 5425, 5427, 5429, 5432, 5434, 5437, 5439, 5442, 5444, 5446, 5449, 5451, 5454, 5456, 5459, 5461, 5464, 5466, 5468, 5471, 5473, 5476, 5478, 5481, 5483, 5486, 5488, 5490, 5493, 5495, 5498, 5500, 5503, 5505, 5508, 5510, 5513, 5515, 5518, 5520, 5522, 5525, 5527, 5530, 5532, 5535, 5537, 5540, 5542, 5545, 5547, 5550, 5552, 5555, 5557, 5560, 5562, 5565, 5567, 5570, 5572, 5575, 5577, 5580, 5582, 5585, 5587, 5590, 5592, 5595, 5597, 5600, 5602, 5605, 5607, 5610, 5612, 5615, 5617, 5620, 5622, 5625, 5627, 5630, 5632, 5635, 5637, 5640, 5642, 5645, 5647, 5650, 5652, 5655, 5657, 5660, 5662, 5665, 5667, 5670, 5672, 5675, 5678, 5680, 5683, 5685, 5688, 5690, 5693, 5695, 5698, 5700, 5703, 5705, 5708, 5711, 5713, 5716, 5718, 5721, 5723, 5726, 5728, 5731, 5733, 5736, 5739, 5741, 5744, 5746, 5749, 5751, 5754, 5757, 5759, 5762, 5764, 5767, 5769, 5772, 5774, 5777, 5780, 5782, 5785, 5787, 5790, 5793, 5795, 5798, 5800, 5803, 5805, 5808, 5811, 5813, 5816, 5818, 5821, 5824, 5826, 5829, 5831, 5834, 5836, 5839, 5842, 5844, 5847, 5849, 5852, 5855, 5857, 5860, 5862, 5865, 5868, 5870, 5873, 5876, 5878, 5881, 5883, 5886, 5889, 5891, 5894, 5896, 5899, 5902, 5904, 5907, 5910, 5912, 5915, 5917, 5920, 5923, 5925, 5928, 5931, 5933, 5936, 5939, 5941, 5944, 5946, 5949, 5952, 5954, 5957, 5960, 5962, 5965, 5968, 5970, 5973, 5976, 5978, 5981, 5984, 5986, 5989, 5991, 5994, 5997, 5999, 6002, 6005, 6007, 6010, 6013, 6015, 6018, 6021, 6023, 6026, 6029, 6031, 6034, 6037, 6039, 6042, 6045, 6048, 6050, 6053, 6056, 6058, 6061, 6064, 6066, 6069, 6072, 6074, 6077, 6080, 6082, 6085, 6088, 6091, 6093, 6096, 6099, 6101, 6104, 6107, 6109, 6112, 6115, 6118, 6120, 6123, 6126, 6128, 6131, 6134, 6137, 6139, 6142, 6145, 6147, 6150, 6153, 6156, 6158, 6161, 6164, 6167, 6169, 6172, 6175, 6177, 6180, 6183, 6186, 6188, 6191, 6194, 6197, 6199, 6202, 6205, 6208, 6210, 6213, 6216, 6219, 6221, 6224, 6227, 6230, 6232, 6235, 6238, 6241, 6243, 6246, 6249, 6252, 6254, 6257, 6260, 6263, 6265, 6268, 6271, 6274, 6276, 6279, 6282, 6285, 6288, 6290, 6293, 6296, 6299, 6301, 6304, 6307, 6310, 6313, 6315, 6318, 6321, 6324, 6327, 6329, 6332, 6335, 6338, 6341, 6343, 6346, 6349, 6352, 6355, 6357, 6360, 6363, 6366, 6369, 6371, 6374, 6377, 6380, 6383, 6385, 6388, 6391, 6394, 6397, 6399, 6402, 6405, 6408, 6411, 6414, 6416, 6419, 6422, 6425, 6428, 6431, 6433, 6436, 6439, 6442, 6445, 6448, 6450, 6453, 6456, 6459, 6462, 6465, 6467, 6470, 6473, 6476, 6479, 6482, 6485, 6487, 6490, 6493, 6496, 6499, 6502, 6505, 6507, 6510, 6513, 6516, 6519, 6522, 6525, 6527, 6530, 6533, 6536, 6539, 6542, 6545, 6548, 6550, 6553, 6556, 6559, 6562, 6565, 6568, 6571, 6574, 6576, 6579, 6582, 6585, 6588, 6591, 6594, 6597, 6600, 6602, 6605, 6608, 6611, 6614, 6617, 6620, 6623, 6626, 6629, 6632, 6634, 6637, 6640, 6643, 6646, 6649, 6652, 6655, 6658, 6661, 6664, 6667, 6669, 6672, 6675, 6678, 6681, 6684, 6687, 6690, 6693, 6696, 6699, 6702, 6705, 6708, 6711, 6713, 6716, 6719, 6722, 6725, 6728, 6731, 6734, 6737, 6740, 6743, 6746, 6749, 6752, 6755, 6758, 6761, 6764, 6767, 6770, 6773, 6776, 6778, 6781, 6784, 6787, 6790, 6793, 6796, 6799, 6802, 6805, 6808, 6811, 6814, 6817, 6820, 6823, 6826, 6829, 6832, 6835, 6838, 6841, 6844, 6847, 6850, 6853, 6856, 6859, 6862, 6865, 6868, 6871, 6874, 6877, 6880, 6883, 6886, 6889, 6892, 6895, 6898, 6901, 6904, 6907, 6910, 6913, 6916, 6919, 6922, 6925, 6928, 6931, 6934, 6937, 6940, 6943, 6946, 6949, 6953, 6956, 6959, 6962, 6965, 6968, 6971, 6974, 6977, 6980, 6983, 6986, 6989, 6992, 6995, 6998, 7001, 7004, 7007, 7010, 7013, 7017, 7020, 7023, 7026, 7029, 7032, 7035, 7038, 7041, 7044, 7047, 7050, 7053, 7056, 7059, 7063, 7066, 7069, 7072, 7075, 7078, 7081, 7084, 7087, 7090, 7093, 7096, 7100, 7103, 7106, 7109, 7112, 7115, 7118, 7121, 7124, 7127, 7131, 7134, 7137, 7140, 7143, 7146, 7149, 7152, 7155, 7158, 7162, 7165, 7168, 7171, 7174, 7177, 7180, 7183, 7187, 7190, 7193, 7196, 7199, 7202, 7205, 7208, 7212, 7215, 7218, 7221, 7224, 7227, 7230, 7234, 7237, 7240, 7243, 7246, 7249, 7252, 7256, 7259, 7262, 7265, 7268, 7271, 7275, 7278, 7281, 7284, 7287, 7290, 7293, 7297, 7300, 7303, 7306, 7309, 7312, 7316, 7319, 7322, 7325, 7328, 7332, 7335, 7338, 7341, 7344, 7347, 7351, 7354, 7357, 7360, 7363, 7367, 7370, 7373, 7376, 7379, 7383, 7386, 7389, 7392, 7395, 7399, 7402, 7405, 7408, 7411, 7415, 7418, 7421, 7424, 7427, 7431, 7434, 7437, 7440, 7444, 7447, 7450, 7453, 7456, 7460, 7463, 7466, 7469, 7473, 7476, 7479, 7482, 7486, 7489, 7492, 7495, 7498, 7502, 7505, 7508, 7511, 7515, 7518, 7521, 7524, 7528, 7531, 7534, 7537, 7541, 7544, 7547, 7551, 7554, 7557, 7560, 7564, 7567, 7570, 7573, 7577, 7580, 7583, 7586, 7590, 7593, 7596, 7600, 7603, 7606, 7609, 7613, 7616, 7619, 7623, 7626, 7629, 7632, 7636, 7639, 7642, 7646, 7649, 7652, 7656, 7659, 7662, 7665, 7669, 7672, 7675, 7679, 7682, 7685, 7689, 7692, 7695, 7699, 7702, 7705, 7709, 7712, 7715, 7718, 7722, 7725, 7728, 7732, 7735, 7738, 7742, 7745, 7748, 7752, 7755, 7758, 7762, 7765, 7769, 7772, 7775, 7779, 7782, 7785, 7789, 7792, 7795, 7799, 7802, 7805, 7809, 7812, 7815, 7819, 7822, 7826, 7829, 7832, 7836, 7839, 7842, 7846, 7849, 7852, 7856, 7859, 7863, 7866, 7869, 7873, 7876, 7880, 7883, 7886, 7890, 7893, 7896, 7900, 7903, 7907, 7910, 7913, 7917, 7920, 7924, 7927, 7930, 7934, 7937, 7941, 7944, 7947, 7951, 7954, 7958, 7961, 7965, 7968, 7971, 7975, 7978, 7982, 7985, 7988, 7992, 7995, 7999, 8002, 8006, 8009, 8012, 8016, 8019, 8023, 8026, 8030, 8033, 8037, 8040, 8043, 8047, 8050, 8054, 8057, 8061, 8064, 8068, 8071, 8075, 8078, 8081, 8085, 8088, 8092, 8095, 8099, 8102, 8106, 8109, 8113, 8116, 8120, 8123, 8127, 8130, 8133, 8137, 8140, 8144, 8147, 8151, 8154, 8158, 8161, 8165, 8168, 8172, 8175, 8179, 8182, 8186, 8189, 8193, 8196, 8200, 8203, 8207, 8210, 8214, 8217, 8221, 8224, 8228, 8231, 8235, 8238, 8242, 8245, 8249, 8252, 8256, 8260, 8263, 8267, 8270, 8274, 8277, 8281, 8284, 8288, 8291, 8295, 8298, 8302, 8305, 8309, 8313, 8316, 8320, 8323, 8327, 8330, 8334, 8337, 8341, 8344, 8348, 8352, 8355, 8359, 8362, 8366, 8369, 8373, 8377, 8380, 8384, 8387, 8391, 8394, 8398, 8402, 8405, 8409, 8412, 8416, 8419, 8423, 8427, 8430, 8434, 8437, 8441, 8445, 8448, 8452, 8455, 8459, 8463, 8466, 8470, 8473, 8477, 8481, 8484, 8488, 8491, 8495, 8499, 8502, 8506, 8509, 8513, 8517, 8520, 8524, 8528, 8531, 8535, 8538, 8542, 8546, 8549, 8553, 8557, 8560, 8564, 8567, 8571, 8575, 8578, 8582, 8586, 8589, 8593, 8597, 8600, 8604, 8608, 8611, 8615, 8618, 8622, 8626, 8629, 8633, 8637, 8640, 8644, 8648, 8651, 8655, 8659, 8662, 8666, 8670, 8673, 8677, 8681, 8684, 8688, 8692, 8696, 8699, 8703, 8707, 8710, 8714, 8718, 8721, 8725, 8729, 8732, 8736, 8740, 8743, 8747, 8751, 8755, 8758, 8762, 8766, 8769, 8773, 8777, 8781, 8784, 8788, 8792, 8795, 8799, 8803, 8807, 8810, 8814, 8818, 8821, 8825, 8829, 8833, 8836, 8840, 8844, 8848, 8851, 8855, 8859, 8863, 8866, 8870, 8874, 8878, 8881, 8885, 8889, 8893, 8896, 8900, 8904, 8908, 8911, 8915, 8919, 8923, 8926, 8930, 8934, 8938, 8941, 8945, 8949, 8953, 8957, 8960, 8964, 8968, 8972, 8975, 8979, 8983, 8987, 8991, 8994, 8998, 9002, 9006, 9010, 9013, 9017, 9021, 9025, 9029, 9032, 9036, 9040, 9044, 9048, 9051, 9055, 9059, 9063, 9067, 9070, 9074, 9078, 9082, 9086, 9090, 9093, 9097, 9101, 9105, 9109, 9112, 9116, 9120, 9124, 9128, 9132, 9135, 9139, 9143, 9147, 9151, 9155, 9159, 9162, 9166, 9170, 9174, 9178, 9182, 9186, 9189, 9193, 9197, 9201, 9205, 9209, 9213, 9216, 9220, 9224, 9228, 9232, 9236, 9240, 9244, 9247, 9251, 9255, 9259, 9263, 9267, 9271, 9275, 9278, 9282, 9286, 9290, 9294, 9298, 9302, 9306, 9310, 9314, 9317, 9321, 9325, 9329, 9333, 9337, 9341, 9345, 9349, 9353, 9357, 9360, 9364, 9368, 9372, 9376, 9380, 9384, 9388, 9392, 9396, 9400, 9404, 9408, 9411, 9415, 9419, 9423, 9427, 9431, 9435, 9439, 9443, 9447, 9451, 9455, 9459, 9463, 9467, 9471, 9475, 9479, 9483, 9486, 9490, 9494, 9498, 9502, 9506, 9510, 9514, 9518, 9522, 9526, 9530, 9534, 9538, 9542, 9546, 9550, 9554, 9558, 9562, 9566, 9570, 9574, 9578, 9582, 9586, 9590, 9594, 9598, 9602, 9606, 9610, 9614, 9618, 9622, 9626, 9630, 9634, 9638, 9642, 9646, 9650, 9654, 9658, 9662, 9666, 9670, 9674, 9678, 9682, 9686, 9690, 9694, 9698, 9702, 9706, 9710, 9715, 9719, 9723, 9727, 9731, 9735, 9739, 9743, 9747, 9751, 9755, 9759, 9763, 9767, 9771, 9775, 9779, 9783, 9787, 9792, 9796, 9800, 9804, 9808, 9812, 9816, 9820, 9824, 9828, 9832, 9836, 9840, 9845, 9849, 9853, 9857, 9861, 9865, 9869, 9873, 9877, 9881, 9885, 9890, 9894, 9898, 9902, 9906, 9910, 9914, 9918, 9922, 9927, 9931, 9935, 9939, 9943, 9947, 9951, 9955, 9959, 9964, 9968, 9972, 9976, 9980, 9984, 9988, 9992, 9997, 10001, 10005, 10009, 10013, 10017, 10021, 10026, 10030, 10034, 10038, 10042, 10046, 10051, 10055, 10059, 10063, 10067, 10071, 10075, 10080, 10084, 10088, 10092, 10096, 10100, 10105, 10109, 10113, 10117, 10121, 10126, 10130, 10134, 10138, 10142, 10146, 10151, 10155, 10159, 10163, 10167, 10172, 10176, 10180, 10184, 10188, 10193, 10197, 10201, 10205, 10209, 10214, 10218, 10222, 10226, 10230, 10235, 10239, 10243, 10247, 10252, 10256, 10260, 10264, 10268, 10273, 10277, 10281, 10285, 10290, 10294, 10298, 10302, 10307, 10311, 10315, 10319, 10324, 10328, 10332, 10336, 10341, 10345, 10349, 10353, 10358, 10362, 10366, 10370, 10375, 10379, 10383, 10387, 10392, 10396, 10400, 10405, 10409, 10413, 10417, 10422, 10426, 10430, 10434, 10439, 10443, 10447, 10452, 10456, 10460, 10464, 10469, 10473, 10477, 10482, 10486, 10490, 10495, 10499, 10503, 10508, 10512, 10516, 10520, 10525, 10529, 10533, 10538, 10542, 10546, 10551, 10555, 10559, 10564, 10568, 10572, 10577, 10581, 10585, 10590, 10594, 10598, 10603, 10607, 10611, 10616, 10620, 10624, 10629, 10633, 10637, 10642, 10646, 10650, 10655, 10659, 10664, 10668, 10672, 10677, 10681, 10685, 10690, 10694, 10698, 10703, 10707, 10712, 10716, 10720, 10725, 10729, 10733, 10738, 10742, 10747, 10751, 10755, 10760, 10764, 10769, 10773, 10777, 10782, 10786, 10791, 10795, 10799, 10804, 10808, 10813, 10817, 10821, 10826, 10830, 10835, 10839, 10843, 10848, 10852, 10857, 10861, 10866, 10870, 10874, 10879, 10883, 10888, 10892, 10897, 10901, 10905, 10910, 10914, 10919, 10923, 10928, 10932, 10937, 10941, 10945, 10950, 10954, 10959, 10963, 10968, 10972, 10977, 10981, 10986, 10990, 10995, 10999, 11003, 11008, 11012, 11017, 11021, 11026, 11030, 11035, 11039, 11044, 11048, 11053, 11057, 11062, 11066, 11071, 11075, 11080, 11084, 11089, 11093, 11098, 11102, 11107, 11111, 11116, 11120, 11125, 11129, 11134, 11138, 11143, 11147, 11152, 11156, 11161, 11165, 11170, 11174, 11179, 11183, 11188, 11193, 11197, 11202, 11206, 11211, 11215, 11220, 11224, 11229, 11233, 11238, 11242, 11247, 11252, 11256, 11261, 11265, 11270, 11274, 11279, 11283, 11288, 11293, 11297, 11302, 11306, 11311, 11315, 11320, 11325, 11329, 11334, 11338, 11343, 11347, 11352, 11357, 11361, 11366, 11370, 11375, 11380, 11384, 11389, 11393, 11398, 11403, 11407, 11412, 11416, 11421, 11426, 11430, 11435, 11439, 11444, 11449, 11453, 11458, 11462, 11467, 11472, 11476, 11481, 11486, 11490, 11495, 11499, 11504, 11509, 11513, 11518, 11523, 11527, 11532, 11537, 11541, 11546, 11550, 11555, 11560, 11564, 11569, 11574, 11578, 11583, 11588, 11592, 11597, 11602, 11606, 11611, 11616, 11620, 11625, 11630, 11634, 11639, 11644, 11648, 11653, 11658, 11662, 11667, 11672, 11676, 11681, 11686, 11690, 11695, 11700, 11705, 11709, 11714, 11719, 11723, 11728, 11733, 11737, 11742, 11747, 11752, 11756, 11761, 11766, 11770, 11775, 11780, 11785, 11789, 11794, 11799, 11803, 11808, 11813, 11818, 11822, 11827, 11832, 11837, 11841, 11846, 11851, 11856, 11860, 11865, 11870, 11875, 11879, 11884, 11889, 11894, 11898, 11903, 11908, 11913, 11917, 11922, 11927, 11932, 11936, 11941, 11946, 11951, 11955, 11960, 11965, 11970, 11975, 11979, 11984, 11989, 11994, 11998, 12003, 12008, 12013, 12018, 12022, 12027, 12032, 12037, 12042, 12046, 12051, 12056, 12061, 12066, 12070, 12075, 12080, 12085, 12090, 12094, 12099, 12104, 12109, 12114, 12119, 12123, 12128, 12133, 12138, 12143, 12148, 12152, 12157, 12162, 12167, 12172, 12177, 12181, 12186, 12191, 12196, 12201, 12206, 12210, 12215, 12220, 12225, 12230, 12235, 12240, 12244, 12249, 12254, 12259, 12264, 12269, 12274, 12279, 12283, 12288, 12293, 12298, 12303, 12308, 12313, 12318, 12322, 12327, 12332, 12337, 12342, 12347, 12352, 12357, 12362, 12366, 12371, 12376, 12381, 12386, 12391, 12396, 12401, 12406, 12411, 12416, 12420, 12425, 12430, 12435, 12440, 12445, 12450, 12455, 12460, 12465, 12470, 12475, 12480, 12484, 12489, 12494, 12499, 12504, 12509, 12514, 12519, 12524, 12529, 12534, 12539, 12544, 12549, 12554, 12559, 12564, 12569, 12574, 12579, 12583, 12588, 12593, 12598, 12603, 12608, 12613, 12618, 12623, 12628, 12633, 12638, 12643, 12648, 12653, 12658, 12663, 12668, 12673, 12678, 12683, 12688, 12693, 12698, 12703, 12708, 12713, 12718, 12723, 12728, 12733, 12738, 12743, 12748, 12753, 12758, 12763, 12768, 12773, 12778, 12783, 12788, 12793, 12798, 12803, 12808, 12813, 12818, 12823, 12829, 12834, 12839, 12844, 12849, 12854, 12859, 12864, 12869, 12874, 12879, 12884, 12889, 12894, 12899, 12904, 12909, 12914, 12919, 12925, 12930, 12935, 12940, 12945, 12950, 12955, 12960, 12965, 12970, 12975, 12980, 12985, 12991, 12996, 13001, 13006, 13011, 13016, 13021, 13026, 13031, 13036, 13041, 13047, 13052, 13057, 13062, 13067, 13072, 13077, 13082, 13087, 13093, 13098, 13103, 13108, 13113, 13118, 13123, 13128, 13133, 13139, 13144, 13149, 13154, 13159, 13164, 13169, 13175, 13180, 13185, 13190, 13195, 13200, 13205, 13211, 13216, 13221, 13226, 13231, 13236, 13242, 13247, 13252, 13257, 13262, 13267, 13272, 13278, 13283, 13288, 13293, 13298, 13304, 13309, 13314, 13319, 13324, 13329, 13335, 13340, 13345, 13350, 13355, 13361, 13366, 13371, 13376, 13381, 13387, 13392, 13397, 13402, 13407, 13413, 13418, 13423, 13428, 13433, 13439, 13444, 13449, 13454, 13460, 13465, 13470, 13475, 13480, 13486, 13491, 13496, 13501, 13507, 13512, 13517, 13522, 13528, 13533, 13538, 13543, 13549, 13554, 13559, 13564, 13570, 13575, 13580, 13585, 13591, 13596, 13601, 13606, 13612, 13617, 13622, 13627, 13633, 13638, 13643, 13648, 13654, 13659, 13664, 13670, 13675, 13680, 13685, 13691, 13696, 13701, 13707, 13712, 13717, 13723, 13728, 13733, 13738, 13744, 13749, 13754, 13760, 13765, 13770, 13776, 13781, 13786, 13792, 13797, 13802, 13807, 13813, 13818, 13823, 13829, 13834, 13839, 13845, 13850, 13855, 13861, 13866, 13871, 13877, 13882, 13887, 13893, 13898, 13903, 13909, 13914, 13920, 13925, 13930, 13936, 13941, 13946, 13952, 13957, 13962, 13968, 13973, 13979, 13984, 13989, 13995, 14000, 14005, 14011, 14016, 14022, 14027, 14032, 14038, 14043, 14048, 14054, 14059, 14065, 14070, 14075, 14081, 14086, 14092, 14097, 14102, 14108, 14113, 14119, 14124, 14129, 14135, 14140, 14146, 14151, 14157, 14162, 14167, 14173, 14178, 14184, 14189, 14195, 14200, 14205, 14211, 14216, 14222, 14227, 14233, 14238, 14243, 14249, 14254, 14260, 14265, 14271, 14276, 14282, 14287, 14292, 14298, 14303, 14309, 14314, 14320, 14325, 14331, 14336, 14342, 14347, 14353, 14358, 14364, 14369, 14375, 14380, 14385, 14391, 14396, 14402, 14407, 14413, 14418, 14424, 14429, 14435, 14440, 14446, 14451, 14457, 14462, 14468, 14473, 14479, 14484, 14490, 14495, 14501, 14506, 14512, 14517, 14523, 14529, 14534, 14540, 14545, 14551, 14556, 14562, 14567, 14573, 14578, 14584, 14589, 14595, 14600, 14606, 14612, 14617, 14623, 14628, 14634, 14639, 14645, 14650, 14656, 14661, 14667, 14673, 14678, 14684, 14689, 14695, 14700, 14706, 14712, 14717, 14723, 14728, 14734, 14739, 14745, 14751, 14756, 14762, 14767, 14773, 14778, 14784, 14790, 14795, 14801, 14806, 14812, 14818, 14823, 14829, 14834, 14840, 14846, 14851, 14857, 14862, 14868, 14874, 14879, 14885, 14891, 14896, 14902, 14907, 14913, 14919, 14924, 14930, 14936, 14941, 14947, 14952, 14958, 14964, 14969, 14975, 14981, 14986, 14992, 14998, 15003, 15009, 15015, 15020, 15026, 15032, 15037, 15043, 15048, 15054, 15060, 15065, 15071, 15077, 15082, 15088, 15094, 15099, 15105, 15111, 15117, 15122, 15128, 15134, 15139, 15145, 15151, 15156, 15162, 15168, 15173, 15179, 15185, 15190, 15196, 15202, 15208, 15213, 15219, 15225, 15230, 15236, 15242, 15248, 15253, 15259, 15265, 15270, 15276, 15282, 15288, 15293, 15299, 15305, 15310, 15316, 15322, 15328, 15333, 15339, 15345, 15351, 15356, 15362, 15368, 15374, 15379, 15385, 15391, 15397, 15402, 15408, 15414, 15420, 15425, 15431, 15437, 15443, 15448, 15454, 15460, 15466, 15471, 15477, 15483, 15489, 15495, 15500, 15506, 15512, 15518, 15523, 15529, 15535, 15541, 15547, 15552, 15558, 15564, 15570, 15576, 15581, 15587, 15593, 15599, 15605, 15610, 15616, 15622, 15628, 15634, 15639, 15645, 15651, 15657, 15663, 15669, 15674, 15680, 15686, 15692, 15698, 15703, 15709, 15715, 15721, 15727, 15733, 15738, 15744, 15750, 15756, 15762, 15768, 15774, 15779, 15785, 15791, 15797, 15803, 15809, 15815, 15820, 15826, 15832, 15838, 15844, 15850, 15856, 15861, 15867, 15873, 15879, 15885, 15891, 15897, 15903, 15908, 15914, 15920, 15926, 15932, 15938, 15944, 15950, 15956, 15961, 15967, 15973, 15979, 15985, 15991, 15997, 16003, 16009, 16015, 16020, 16026, 16032, 16038, 16044, 16050, 16056, 16062, 16068, 16074, 16080, 16086, 16092, 16097, 16103, 16109, 16115, 16121, 16127, 16133, 16139, 16145, 16151, 16157, 16163, 16169, 16175, 16181, 16187, 16193, 16198, 16204, 16210, 16216, 16222, 16228, 16234, 16240, 16246, 16252, 16258, 16264, 16270, 16276, 16282, 16288, 16294, 16300, 16306, 16312, 16318, 16324, 16330, 16336, 16342, 16348, 16354, 16360, 16366, 16372, 16378, 16384, 16390, 16396, 16402, 16408, 16414, 16420, 16426, 16432, 16438, 16444, 16450, 16456, 16462, 16468, 16474, 16480, 16486, 16492, 16498, 16504, 16510, 16516, 16522, 16528, 16534, 16540, 16546, 16552, 16558, 16564, 16570, 16576, 16583, 16589, 16595, 16601, 16607, 16613, 16619, 16625, 16631, 16637, 16643, 16649, 16655, 16661, 16667, 16673, 16679, 16686, 16692, 16698, 16704, 16710, 16716, 16722, 16728, 16734, 16740, 16746, 16752, 16759, 16765, 16771, 16777, 16783, 16789, 16795, 16801, 16807, 16813, 16820, 16826, 16832, 16838, 16844, 16850, 16856, 16862, 16868, 16875, 16881, 16887, 16893, 16899, 16905, 16911, 16917, 16924, 16930, 16936, 16942, 16948, 16954, 16960, 16966, 16973, 16979, 16985, 16991, 16997, 17003, 17009, 17016, 17022, 17028, 17034, 17040, 17046, 17053, 17059, 17065, 17071, 17077, 17083, 17090, 17096, 17102, 17108, 17114, 17120, 17127, 17133, 17139, 17145, 17151, 17157, 17164, 17170, 17176, 17182, 17188, 17195, 17201, 17207, 17213, 17219, 17226, 17232, 17238, 17244, 17250, 17257, 17263, 17269, 17275, 17281, 17288, 17294, 17300, 17306, 17313, 17319, 17325, 17331, 17337, 17344, 17350, 17356, 17362, 17369, 17375, 17381, 17387, 17394, 17400, 17406, 17412, 17418, 17425, 17431, 17437, 17443, 17450, 17456, 17462, 17468, 17475, 17481, 17487, 17494, 17500, 17506, 17512, 17519, 17525, 17531, 17537, 17544, 17550, 17556, 17563, 17569, 17575, 17581, 17588, 17594, 17600, 17606, 17613, 17619, 17625, 17632, 17638, 17644, 17651, 17657, 17663, 17669, 17676, 17682, 17688, 17695, 17701, 17707, 17714, 17720, 17726, 17733, 17739, 17745, 17751, 17758, 17764, 17770, 17777, 17783, 17789, 17796, 17802, 17808, 17815, 17821, 17827, 17834, 17840, 17846, 17853, 17859, 17865, 17872, 17878, 17884, 17891, 17897, 17904, 17910, 17916, 17923, 17929, 17935, 17942, 17948, 17954, 17961, 17967, 17974, 17980, 17986, 17993, 17999, 18005, 18012, 18018, 18025, 18031, 18037, 18044, 18050, 18056, 18063, 18069, 18076, 18082, 18088, 18095, 18101, 18108, 18114, 18120, 18127, 18133, 18140, 18146, 18152, 18159, 18165, 18172, 18178, 18184, 18191, 18197, 18204, 18210, 18217, 18223, 18229, 18236, 18242, 18249, 18255, 18262, 18268, 18274, 18281, 18287, 18294, 18300, 18307, 18313, 18319, 18326, 18332, 18339, 18345, 18352, 18358, 18365, 18371, 18378, 18384, 18390, 18397, 18403, 18410, 18416, 18423, 18429, 18436, 18442, 18449, 18455, 18462, 18468, 18475, 18481, 18488, 18494, 18500, 18507, 18513, 18520, 18526, 18533, 18539, 18546, 18552, 18559, 18565, 18572, 18578, 18585, 18591, 18598, 18604, 18611, 18617, 18624, 18630, 18637, 18643, 18650, 18656, 18663, 18670, 18676, 18683, 18689, 18696, 18702, 18709, 18715, 18722, 18728, 18735, 18741, 18748, 18754, 18761, 18767, 18774, 18781, 18787, 18794, 18800, 18807, 18813, 18820, 18826, 18833, 18839, 18846, 18853, 18859, 18866, 18872, 18879, 18885, 18892, 18899, 18905, 18912, 18918, 18925, 18931, 18938, 18945, 18951, 18958, 18964, 18971, 18977, 18984, 18991, 18997, 19004, 19010, 19017, 19024, 19030, 19037, 19043, 19050, 19057, 19063, 19070, 19076, 19083, 19090, 19096, 19103, 19109, 19116, 19123, 19129, 19136, 19142, 19149, 19156, 19162, 19169, 19176, 19182, 19189, 19195, 19202, 19209, 19215, 19222, 19229, 19235, 19242, 19248, 19255, 19262, 19268, 19275, 19282, 19288, 19295, 19302, 19308, 19315, 19322, 19328, 19335, 19342, 19348, 19355, 19362, 19368, 19375, 19381, 19388, 19395, 19401, 19408, 19415, 19422, 19428, 19435, 19442, 19448, 19455, 19462, 19468, 19475, 19482, 19488, 19495, 19502, 19508, 19515, 19522, 19528, 19535, 19542, 19549, 19555, 19562, 19569, 19575, 19582, 19589, 19595, 19602, 19609, 19616, 19622, 19629, 19636, 19642, 19649, 19656, 19663, 19669, 19676, 19683, 19689, 19696, 19703, 19710, 19716, 19723, 19730, 19737, 19743, 19750, 19757, 19764, 19770, 19777, 19784, 19791, 19797, 19804, 19811, 19818, 19824, 19831, 19838, 19845, 19851, 19858, 19865, 19872, 19878, 19885, 19892, 19899, 19905, 19912, 19919, 19926, 19932, 19939, 19946, 19953, 19960, 19966, 19973, 19980, 19987, 19993, 20000, 20007, 20014, 20021, 20027, 20034, 20041, 20048, 20055, 20061, 20068, 20075, 20082, 20089, 20095, 20102, 20109, 20116, 20123, 20129, 20136, 20143, 20150, 20157, 20163, 20170, 20177, 20184, 20191, 20198, 20204, 20211, 20218, 20225, 20232, 20239, 20245, 20252, 20259, 20266, 20273, 20280, 20286, 20293, 20300, 20307, 20314, 20321, 20327, 20334, 20341, 20348, 20355, 20362, 20369, 20375, 20382, 20389, 20396, 20403, 20410, 20417, 20423, 20430, 20437, 20444, 20451, 20458, 20465, 20471, 20478, 20485, 20492, 20499, 20506, 20513, 20520, 20527, 20533, 20540, 20547, 20554, 20561, 20568, 20575, 20582, 20589, 20595, 20602, 20609, 20616, 20623, 20630, 20637, 20644, 20651, 20658, 20664, 20671, 20678, 20685, 20692, 20699, 20706, 20713, 20720, 20727, 20734, 20740, 20747, 20754, 20761, 20768, 20775, 20782, 20789, 20796, 20803, 20810, 20817, 20824, 20831, 20838, 20844, 20851, 20858, 20865, 20872, 20879, 20886, 20893, 20900, 20907, 20914, 20921, 20928, 20935, 20942, 20949, 20956, 20963, 20970, 20977, 20984, 20990, 20997, 21004, 21011, 21018, 21025, 21032, 21039, 21046, 21053, 21060, 21067, 21074, 21081, 21088, 21095, 21102, 21109, 21116, 21123, 21130, 21137, 21144, 21151, 21158, 21165, 21172, 21179, 21186, 21193, 21200, 21207, 21214, 21221, 21228, 21235, 21242, 21249, 21256, 21263, 21270, 21277, 21284, 21291, 21298, 21305, 21312, 21319, 21326, 21333, 21340, 21347, 21354, 21361, 21368, 21375, 21383, 21390, 21397, 21404, 21411, 21418, 21425, 21432, 21439, 21446, 21453, 21460, 21467, 21474, 21481, 21488, 21495, 21502, 21509, 21516, 21523, 21531, 21538, 21545, 21552, 21559, 21566, 21573, 21580, 21587, 21594, 21601, 21608, 21615, 21622, 21629, 21637, 21644, 21651, 21658, 21665, 21672, 21679, 21686, 21693, 21700, 21707, 21714, 21722, 21729, 21736, 21743, 21750, 21757, 21764, 21771, 21778, 21785, 21792, 21800, 21807, 21814, 21821, 21828, 21835, 21842, 21849, 21856, 21864, 21871, 21878, 21885, 21892, 21899, 21906, 21913, 21921, 21928, 21935, 21942, 21949, 21956, 21963, 21970, 21978, 21985, 21992, 21999, 22006, 22013, 22020, 22028, 22035, 22042, 22049, 22056, 22063, 22070, 22078, 22085, 22092, 22099, 22106, 22113, 22120, 22128, 22135, 22142, 22149, 22156, 22163, 22171, 22178, 22185, 22192, 22199, 22206, 22214, 22221, 22228, 22235, 22242, 22249, 22257, 22264, 22271, 22278, 22285, 22292, 22300, 22307, 22314, 22321, 22328, 22336, 22343, 22350, 22357, 22364, 22372, 22379, 22386, 22393, 22400, 22408, 22415, 22422, 22429, 22436, 22444, 22451, 22458, 22465, 22472, 22480, 22487, 22494, 22501, 22508, 22516, 22523, 22530, 22537, 22545, 22552, 22559, 22566, 22573, 22581, 22588, 22595, 22602, 22610, 22617, 22624, 22631, 22639, 22646, 22653, 22660, 22667, 22675, 22682, 22689, 22696, 22704, 22711, 22718, 22725, 22733, 22740, 22747, 22754, 22762, 22769, 22776, 22783, 22791, 22798, 22805, 22812, 22820, 22827, 22834, 22842, 22849, 22856, 22863, 22871, 22878, 22885, 22892, 22900, 22907, 22914, 22922, 22929, 22936, 22943, 22951, 22958, 22965, 22973, 22980, 22987, 22994, 23002, 23009, 23016, 23024, 23031, 23038, 23045, 23053, 23060, 23067, 23075, 23082, 23089, 23097, 23104, 23111, 23118, 23126, 23133, 23140, 23148, 23155, 23162, 23170, 23177, 23184, 23192, 23199, 23206, 23213, 23221, 23228, 23235, 23243, 23250, 23257, 23265, 23272, 23279, 23287, 23294, 23301, 23309, 23316, 23323, 23331, 23338, 23345, 23353, 23360, 23367, 23375, 23382, 23389, 23397, 23404, 23411, 23419, 23426, 23434, 23441, 23448, 23456, 23463, 23470, 23478, 23485, 23492, 23500, 23507, 23514, 23522, 23529, 23537, 23544, 23551, 23559, 23566, 23573, 23581, 23588, 23596, 23603, 23610, 23618, 23625, 23632, 23640, 23647, 23655, 23662, 23669, 23677, 23684, 23691, 23699, 23706, 23714, 23721, 23728, 23736, 23743, 23751, 23758, 23765, 23773, 23780, 23788, 23795, 23802, 23810, 23817, 23825, 23832, 23839, 23847, 23854, 23862, 23869, 23876, 23884, 23891, 23899, 23906, 23913, 23921, 23928, 23936, 23943, 23951, 23958, 23965, 23973, 23980, 23988, 23995, 24003, 24010, 24017, 24025, 24032, 24040, 24047, 24055, 24062, 24069, 24077, 24084, 24092, 24099, 24107, 24114, 24122, 24129, 24136, 24144, 24151, 24159, 24166, 24174, 24181, 24189, 24196, 24203, 24211, 24218, 24226, 24233, 24241, 24248, 24256, 24263, 24271, 24278, 24285, 24293, 24300, 24308, 24315, 24323, 24330, 24338, 24345, 24353, 24360, 24368, 24375, 24383, 24390, 24398, 24405, 24413, 24420, 24427, 24435, 24442, 24450, 24457, 24465, 24472, 24480, 24487, 24495, 24502, 24510, 24517, 24525, 24532, 24540, 24547, 24555, 24562, 24570, 24577, 24585, 24592, 24600, 24607, 24615, 24622, 24630, 24637, 24645, 24652, 24660, 24667, 24675, 24682, 24690, 24697, 24705, 24712, 24720, 24727, 24735, 24743, 24750, 24758, 24765, 24773, 24780, 24788, 24795, 24803, 24810, 24818, 24825, 24833, 24840, 24848, 24855, 24863, 24870, 24878, 24886, 24893, 24901, 24908, 24916, 24923, 24931, 24938, 24946, 24953, 24961, 24969, 24976, 24984, 24991, 24999, 25006, 25014, 25021, 25029, 25036, 25044, 25052, 25059, 25067, 25074, 25082, 25089, 25097, 25104, 25112, 25120, 25127, 25135, 25142, 25150, 25157, 25165, 25173, 25180, 25188, 25195, 25203, 25210, 25218, 25226, 25233, 25241, 25248, 25256, 25263, 25271, 25279, 25286, 25294, 25301, 25309, 25317, 25324, 25332, 25339, 25347, 25355, 25362, 25370, 25377, 25385, 25392, 25400, 25408, 25415, 25423, 25430, 25438, 25446, 25453, 25461, 25468, 25476, 25484, 25491, 25499, 25506, 25514, 25522, 25529, 25537, 25545, 25552, 25560, 25567, 25575, 25583, 25590, 25598, 25605, 25613, 25621, 25628, 25636, 25644, 25651, 25659, 25666, 25674, 25682, 25689, 25697, 25705, 25712, 25720, 25727, 25735, 25743, 25750, 25758, 25766, 25773, 25781, 25789, 25796, 25804, 25811, 25819, 25827, 25834, 25842, 25850, 25857, 25865, 25873, 25880, 25888, 25896, 25903, 25911, 25918, 25926, 25934, 25941, 25949, 25957, 25964, 25972, 25980, 25987, 25995, 26003, 26010, 26018, 26026, 26033, 26041, 26049, 26056, 26064, 26072, 26079, 26087, 26095, 26102, 26110, 26118, 26125, 26133, 26141, 26148, 26156, 26164, 26171, 26179, 26187, 26194, 26202, 26210, 26217, 26225, 26233, 26240, 26248, 26256, 26264, 26271, 26279, 26287, 26294, 26302, 26310, 26317, 26325, 26333, 26340, 26348, 26356, 26363, 26371, 26379, 26387, 26394, 26402, 26410, 26417, 26425, 26433, 26440, 26448, 26456, 26464, 26471, 26479, 26487, 26494, 26502, 26510, 26518, 26525, 26533, 26541, 26548, 26556, 26564, 26571, 26579, 26587, 26595, 26602, 26610, 26618, 26626, 26633, 26641, 26649, 26656, 26664, 26672, 26680, 26687, 26695, 26703, 26710, 26718, 26726, 26734, 26741, 26749, 26757, 26765, 26772, 26780, 26788, 26795, 26803, 26811, 26819, 26826, 26834, 26842, 26850, 26857, 26865, 26873, 26881, 26888, 26896, 26904, 26912, 26919, 26927, 26935, 26943, 26950, 26958, 26966, 26974, 26981, 26989, 26997, 27005, 27012, 27020, 27028, 27036, 27043, 27051, 27059, 27067, 27074, 27082, 27090, 27098, 27105, 27113, 27121, 27129, 27136, 27144, 27152, 27160, 27168, 27175, 27183, 27191, 27199, 27206, 27214, 27222, 27230, 27237, 27245, 27253, 27261, 27269, 27276, 27284, 27292, 27300, 27307, 27315, 27323, 27331, 27339, 27346, 27354, 27362, 27370, 27377, 27385, 27393, 27401, 27409, 27416, 27424, 27432, 27440, 27448, 27455, 27463, 27471, 27479, 27486, 27494, 27502, 27510, 27518, 27525, 27533, 27541, 27549, 27557, 27564, 27572, 27580, 27588, 27596, 27603, 27611, 27619, 27627, 27635, 27642, 27650, 27658, 27666, 27674, 27681, 27689, 27697, 27705, 27713, 27720, 27728, 27736, 27744, 27752, 27760, 27767, 27775, 27783, 27791, 27799, 27806, 27814, 27822, 27830, 27838, 27846, 27853, 27861, 27869, 27877, 27885, 27892, 27900, 27908, 27916, 27924, 27932, 27939, 27947, 27955, 27963, 27971, 27979, 27986, 27994, 28002, 28010, 28018, 28026, 28033, 28041, 28049, 28057, 28065, 28073, 28080, 28088, 28096, 28104, 28112, 28120, 28127, 28135, 28143, 28151, 28159, 28167, 28174, 28182, 28190, 28198, 28206, 28214, 28222, 28229, 28237, 28245, 28253, 28261, 28269, 28276, 28284, 28292, 28300, 28308, 28316, 28324, 28331, 28339, 28347, 28355, 28363, 28371, 28379, 28386, 28394, 28402, 28410, 28418, 28426, 28434, 28441, 28449, 28457, 28465, 28473, 28481, 28489, 28496, 28504, 28512, 28520, 28528, 28536, 28544, 28552, 28559, 28567, 28575, 28583, 28591, 28599, 28607, 28614, 28622, 28630, 28638, 28646, 28654, 28662, 28670, 28677, 28685, 28693, 28701, 28709, 28717, 28725, 28733, 28740, 28748, 28756, 28764, 28772, 28780, 28788, 28796, 28804, 28811, 28819, 28827, 28835, 28843, 28851, 28859, 28867, 28874, 28882, 28890, 28898, 28906, 28914, 28922, 28930, 28938, 28945, 28953, 28961, 28969, 28977, 28985, 28993, 29001, 29009, 29017, 29024, 29032, 29040, 29048, 29056, 29064, 29072, 29080, 29088, 29095, 29103, 29111, 29119, 29127, 29135, 29143, 29151, 29159, 29167, 29175, 29182, 29190, 29198, 29206, 29214, 29222, 29230, 29238, 29246, 29254, 29261, 29269, 29277, 29285, 29293, 29301, 29309, 29317, 29325, 29333, 29341, 29348, 29356, 29364, 29372, 29380, 29388, 29396, 29404, 29412, 29420, 29428, 29436, 29443, 29451, 29459, 29467, 29475, 29483, 29491, 29499, 29507, 29515, 29523, 29531, 29539, 29546, 29554, 29562, 29570, 29578, 29586, 29594, 29602, 29610, 29618, 29626, 29634, 29642, 29649, 29657, 29665, 29673, 29681, 29689, 29697, 29705, 29713, 29721, 29729, 29737, 29745, 29753, 29760, 29768, 29776, 29784, 29792, 29800, 29808, 29816, 29824, 29832, 29840, 29848, 29856, 29864, 29872, 29880, 29887, 29895, 29903, 29911, 29919, 29927, 29935, 29943, 29951, 29959, 29967, 29975, 29983, 29991, 29999, 30007, 30015, 30022, 30030, 30038, 30046, 30054, 30062, 30070, 30078, 30086, 30094, 30102, 30110, 30118, 30126, 30134, 30142, 30150, 30158, 30165, 30173, 30181, 30189, 30197, 30205, 30213, 30221, 30229, 30237, 30245, 30253, 30261, 30269, 30277, 30285, 30293, 30301, 30309, 30317, 30325, 30332, 30340, 30348, 30356, 30364, 30372, 30380, 30388, 30396, 30404, 30412, 30420, 30428, 30436, 30444, 30452, 30460, 30468, 30476, 30484, 30492, 30500, 30508, 30516, 30524, 30531, 30539, 30547, 30555, 30563, 30571, 30579, 30587, 30595, 30603, 30611, 30619, 30627, 30635, 30643, 30651, 30659, 30667, 30675, 30683, 30691, 30699, 30707, 30715, 30723, 30731, 30739, 30747, 30755, 30763, 30770, 30778, 30786, 30794, 30802, 30810, 30818, 30826, 30834, 30842, 30850, 30858, 30866, 30874, 30882, 30890, 30898, 30906, 30914, 30922, 30930, 30938, 30946, 30954, 30962, 30970, 30978, 30986, 30994, 31002, 31010, 31018, 31026, 31034, 31042, 31050, 31058, 31066, 31074, 31081, 31089, 31097, 31105, 31113, 31121, 31129, 31137, 31145, 31153, 31161, 31169, 31177, 31185, 31193, 31201, 31209, 31217, 31225, 31233, 31241, 31249, 31257, 31265, 31273, 31281, 31289, 31297, 31305, 31313, 31321, 31329, 31337, 31345, 31353, 31361, 31369, 31377, 31385, 31393, 31401, 31409, 31417, 31425, 31433, 31441, 31449, 31457, 31465, 31473, 31481, 31489, 31497, 31505, 31513, 31521, 31529, 31537, 31545, 31553, 31561, 31569, 31577, 31585, 31593, 31600, 31608, 31616, 31624, 31632, 31640, 31648, 31656, 31664, 31672, 31680, 31688, 31696, 31704, 31712, 31720, 31728, 31736, 31744, 31752, 31760, 31768, 31776, 31784, 31792, 31800, 31808, 31816, 31824, 31832, 31840, 31848, 31856, 31864, 31872, 31880, 31888, 31896, 31904, 31912, 31920, 31928, 31936, 31944, 31952, 31960, 31968, 31976, 31984, 31992, 32000, 32008, 32016, 32024, 32032, 32040, 32048, 32056, 32064, 32072, 32080, 32088, 32096, 32104, 32112, 32120, 32128, 32136, 32144, 32152, 32160, 32168, 32176, 32184, 32192, 32200, 32208, 32216, 32224, 32232, 32240, 32248, 32256, 32264, 32272, 32280, 32288, 32296, 32304, 32312, 32320, 32328, 32336, 32344, 32352, 32360, 32368, 32376, 32384, 32392, 32400, 32408, 32416, 32424, 32432, 32440, 32448, 32456, 32464, 32472, 32480, 32488, 32496, 32504, 32512, 32520, 32528, 32536, 32544, 32552, 32560, 32568, 32576, 32584, 32592, 32600, 32608, 32616, 32624, 32632, 32640, 32648, 32656, 32664, 32672, 32680, 32688, 32696, 32704, 32712, 32720, 32728, 32736, 32744, 32752, 32760, 32768, 32776, 32784, 32792, 32800, 32808, 32816, 32824, 32832, 32840, 32848, 32856, 32864, 32872, 32880, 32888, 32896, 32904, 32912, 32920, 32928, 32936, 32944, 32952, 32960, 32968, 32976, 32984, 32992, 33000, 33008, 33016, 33024, 33032, 33040, 33048, 33056, 33064, 33072, 33080, 33088, 33096, 33104, 33112, 33120, 33128, 33136, 33144, 33152, 33160, 33168, 33176, 33184, 33192, 33200, 33208, 33216, 33224, 33232, 33240, 33248, 33256, 33264, 33272, 33280, 33288, 33296, 33304, 33312, 33320, 33328, 33336, 33344, 33352, 33360, 33368, 33376, 33384, 33392, 33400, 33408, 33416, 33424, 33432, 33440, 33448, 33456, 33464, 33472, 33480, 33488, 33496, 33504, 33512, 33520, 33528, 33536, 33544, 33552, 33560, 33568, 33576, 33584, 33592, 33600, 33608, 33616, 33624, 33632, 33640, 33648, 33656, 33664, 33672, 33680, 33688, 33696, 33704, 33712, 33720, 33728, 33736, 33744, 33752, 33760, 33768, 33776, 33784, 33792, 33800, 33808, 33816, 33824, 33832, 33840, 33848, 33856, 33864, 33872, 33880, 33888, 33896, 33904, 33912, 33920, 33928, 33936, 33943, 33951, 33959, 33967, 33975, 33983, 33991, 33999, 34007, 34015, 34023, 34031, 34039, 34047, 34055, 34063, 34071, 34079, 34087, 34095, 34103, 34111, 34119, 34127, 34135, 34143, 34151, 34159, 34167, 34175, 34183, 34191, 34199, 34207, 34215, 34223, 34231, 34239, 34247, 34255, 34263, 34271, 34279, 34287, 34295, 34303, 34311, 34319, 34327, 34335, 34343, 34351, 34359, 34367, 34375, 34383, 34391, 34399, 34407, 34415, 34423, 34431, 34439, 34447, 34455, 34462, 34470, 34478, 34486, 34494, 34502, 34510, 34518, 34526, 34534, 34542, 34550, 34558, 34566, 34574, 34582, 34590, 34598, 34606, 34614, 34622, 34630, 34638, 34646, 34654, 34662, 34670, 34678, 34686, 34694, 34702, 34710, 34718, 34726, 34734, 34742, 34750, 34758, 34766, 34773, 34781, 34789, 34797, 34805, 34813, 34821, 34829, 34837, 34845, 34853, 34861, 34869, 34877, 34885, 34893, 34901, 34909, 34917, 34925, 34933, 34941, 34949, 34957, 34965, 34973, 34981, 34989, 34997, 35005, 35012, 35020, 35028, 35036, 35044, 35052, 35060, 35068, 35076, 35084, 35092, 35100, 35108, 35116, 35124, 35132, 35140, 35148, 35156, 35164, 35172, 35180, 35188, 35196, 35204, 35211, 35219, 35227, 35235, 35243, 35251, 35259, 35267, 35275, 35283, 35291, 35299, 35307, 35315, 35323, 35331, 35339, 35347, 35355, 35363, 35371, 35378, 35386, 35394, 35402, 35410, 35418, 35426, 35434, 35442, 35450, 35458, 35466, 35474, 35482, 35490, 35498, 35506, 35514, 35521, 35529, 35537, 35545, 35553, 35561, 35569, 35577, 35585, 35593, 35601, 35609, 35617, 35625, 35633, 35641, 35649, 35656, 35664, 35672, 35680, 35688, 35696, 35704, 35712, 35720, 35728, 35736, 35744, 35752, 35760, 35768, 35776, 35783, 35791, 35799, 35807, 35815, 35823, 35831, 35839, 35847, 35855, 35863, 35871, 35879, 35887, 35894, 35902, 35910, 35918, 35926, 35934, 35942, 35950, 35958, 35966, 35974, 35982, 35990, 35997, 36005, 36013, 36021, 36029, 36037, 36045, 36053, 36061, 36069, 36077, 36085, 36093, 36100, 36108, 36116, 36124, 36132, 36140, 36148, 36156, 36164, 36172, 36180, 36188, 36195, 36203, 36211, 36219, 36227, 36235, 36243, 36251, 36259, 36267, 36275, 36282, 36290, 36298, 36306, 36314, 36322, 36330, 36338, 36346, 36354, 36361, 36369, 36377, 36385, 36393, 36401, 36409, 36417, 36425, 36433, 36441, 36448, 36456, 36464, 36472, 36480, 36488, 36496, 36504, 36512, 36519, 36527, 36535, 36543, 36551, 36559, 36567, 36575, 36583, 36591, 36598, 36606, 36614, 36622, 36630, 36638, 36646, 36654, 36662, 36669, 36677, 36685, 36693, 36701, 36709, 36717, 36725, 36732, 36740, 36748, 36756, 36764, 36772, 36780, 36788, 36796, 36803, 36811, 36819, 36827, 36835, 36843, 36851, 36859, 36866, 36874, 36882, 36890, 36898, 36906, 36914, 36922, 36929, 36937, 36945, 36953, 36961, 36969, 36977, 36984, 36992, 37000, 37008, 37016, 37024, 37032, 37040, 37047, 37055, 37063, 37071, 37079, 37087, 37095, 37102, 37110, 37118, 37126, 37134, 37142, 37150, 37157, 37165, 37173, 37181, 37189, 37197, 37205, 37212, 37220, 37228, 37236, 37244, 37252, 37260, 37267, 37275, 37283, 37291, 37299, 37307, 37314, 37322, 37330, 37338, 37346, 37354, 37362, 37369, 37377, 37385, 37393, 37401, 37409, 37416, 37424, 37432, 37440, 37448, 37456, 37463, 37471, 37479, 37487, 37495, 37503, 37510, 37518, 37526, 37534, 37542, 37550, 37557, 37565, 37573, 37581, 37589, 37597, 37604, 37612, 37620, 37628, 37636, 37644, 37651, 37659, 37667, 37675, 37683, 37690, 37698, 37706, 37714, 37722, 37730, 37737, 37745, 37753, 37761, 37769, 37776, 37784, 37792, 37800, 37808, 37816, 37823, 37831, 37839, 37847, 37855, 37862, 37870, 37878, 37886, 37894, 37901, 37909, 37917, 37925, 37933, 37940, 37948, 37956, 37964, 37972, 37979, 37987, 37995, 38003, 38011, 38018, 38026, 38034, 38042, 38050, 38057, 38065, 38073, 38081, 38088, 38096, 38104, 38112, 38120, 38127, 38135, 38143, 38151, 38159, 38166, 38174, 38182, 38190, 38197, 38205, 38213, 38221, 38229, 38236, 38244, 38252, 38260, 38267, 38275, 38283, 38291, 38299, 38306, 38314, 38322, 38330, 38337, 38345, 38353, 38361, 38368, 38376, 38384, 38392, 38400, 38407, 38415, 38423, 38431, 38438, 38446, 38454, 38462, 38469, 38477, 38485, 38493, 38500, 38508, 38516, 38524, 38531, 38539, 38547, 38555, 38562, 38570, 38578, 38586, 38593, 38601, 38609, 38617, 38624, 38632, 38640, 38648, 38655, 38663, 38671, 38679, 38686, 38694, 38702, 38710, 38717, 38725, 38733, 38741, 38748, 38756, 38764, 38771, 38779, 38787, 38795, 38802, 38810, 38818, 38826, 38833, 38841, 38849, 38856, 38864, 38872, 38880, 38887, 38895, 38903, 38910, 38918, 38926, 38934, 38941, 38949, 38957, 38965, 38972, 38980, 38988, 38995, 39003, 39011, 39018, 39026, 39034, 39042, 39049, 39057, 39065, 39072, 39080, 39088, 39096, 39103, 39111, 39119, 39126, 39134, 39142, 39149, 39157, 39165, 39173, 39180, 39188, 39196, 39203, 39211, 39219, 39226, 39234, 39242, 39249, 39257, 39265, 39272, 39280, 39288, 39296, 39303, 39311, 39319, 39326, 39334, 39342, 39349, 39357, 39365, 39372, 39380, 39388, 39395, 39403, 39411, 39418, 39426, 39434, 39441, 39449, 39457, 39464, 39472, 39480, 39487, 39495, 39503, 39510, 39518, 39526, 39533, 39541, 39549, 39556, 39564, 39572, 39579, 39587, 39595, 39602, 39610, 39618, 39625, 39633, 39640, 39648, 39656, 39663, 39671, 39679, 39686, 39694, 39702, 39709, 39717, 39725, 39732, 39740, 39747, 39755, 39763, 39770, 39778, 39786, 39793, 39801, 39809, 39816, 39824, 39831, 39839, 39847, 39854, 39862, 39870, 39877, 39885, 39892, 39900, 39908, 39915, 39923, 39931, 39938, 39946, 39953, 39961, 39969, 39976, 39984, 39991, 39999, 40007, 40014, 40022, 40030, 40037, 40045, 40052, 40060, 40068, 40075, 40083, 40090, 40098, 40106, 40113, 40121, 40128, 40136, 40144, 40151, 40159, 40166, 40174, 40181, 40189, 40197, 40204, 40212, 40219, 40227, 40235, 40242, 40250, 40257, 40265, 40273, 40280, 40288, 40295, 40303, 40310, 40318, 40326, 40333, 40341, 40348, 40356, 40363, 40371, 40379, 40386, 40394, 40401, 40409, 40416, 40424, 40432, 40439, 40447, 40454, 40462, 40469, 40477, 40484, 40492, 40500, 40507, 40515, 40522, 40530, 40537, 40545, 40552, 40560, 40567, 40575, 40583, 40590, 40598, 40605, 40613, 40620, 40628, 40635, 40643, 40650, 40658, 40666, 40673, 40681, 40688, 40696, 40703, 40711, 40718, 40726, 40733, 40741, 40748, 40756, 40763, 40771, 40778, 40786, 40793, 40801, 40809, 40816, 40824, 40831, 40839, 40846, 40854, 40861, 40869, 40876, 40884, 40891, 40899, 40906, 40914, 40921, 40929, 40936, 40944, 40951, 40959, 40966, 40974, 40981, 40989, 40996, 41004, 41011, 41019, 41026, 41034, 41041, 41049, 41056, 41064, 41071, 41079, 41086, 41094, 41101, 41109, 41116, 41123, 41131, 41138, 41146, 41153, 41161, 41168, 41176, 41183, 41191, 41198, 41206, 41213, 41221, 41228, 41236, 41243, 41251, 41258, 41265, 41273, 41280, 41288, 41295, 41303, 41310, 41318, 41325, 41333, 41340, 41347, 41355, 41362, 41370, 41377, 41385, 41392, 41400, 41407, 41414, 41422, 41429, 41437, 41444, 41452, 41459, 41467, 41474, 41481, 41489, 41496, 41504, 41511, 41519, 41526, 41533, 41541, 41548, 41556, 41563, 41571, 41578, 41585, 41593, 41600, 41608, 41615, 41623, 41630, 41637, 41645, 41652, 41660, 41667, 41674, 41682, 41689, 41697, 41704, 41711, 41719, 41726, 41734, 41741, 41748, 41756, 41763, 41771, 41778, 41785, 41793, 41800, 41808, 41815, 41822, 41830, 41837, 41845, 41852, 41859, 41867, 41874, 41881, 41889, 41896, 41904, 41911, 41918, 41926, 41933, 41940, 41948, 41955, 41963, 41970, 41977, 41985, 41992, 41999, 42007, 42014, 42022, 42029, 42036, 42044, 42051, 42058, 42066, 42073, 42080, 42088, 42095, 42102, 42110, 42117, 42125, 42132, 42139, 42147, 42154, 42161, 42169, 42176, 42183, 42191, 42198, 42205, 42213, 42220, 42227, 42235, 42242, 42249, 42257, 42264, 42271, 42279, 42286, 42293, 42301, 42308, 42315, 42323, 42330, 42337, 42344, 42352, 42359, 42366, 42374, 42381, 42388, 42396, 42403, 42410, 42418, 42425, 42432, 42439, 42447, 42454, 42461, 42469, 42476, 42483, 42491, 42498, 42505, 42512, 42520, 42527, 42534, 42542, 42549, 42556, 42563, 42571, 42578, 42585, 42593, 42600, 42607, 42614, 42622, 42629, 42636, 42644, 42651, 42658, 42665, 42673, 42680, 42687, 42694, 42702, 42709, 42716, 42724, 42731, 42738, 42745, 42753, 42760, 42767, 42774, 42782, 42789, 42796, 42803, 42811, 42818, 42825, 42832, 42840, 42847, 42854, 42861, 42869, 42876, 42883, 42890, 42897, 42905, 42912, 42919, 42926, 42934, 42941, 42948, 42955, 42963, 42970, 42977, 42984, 42991, 42999, 43006, 43013, 43020, 43028, 43035, 43042, 43049, 43056, 43064, 43071, 43078, 43085, 43092, 43100, 43107, 43114, 43121, 43128, 43136, 43143, 43150, 43157, 43164, 43172, 43179, 43186, 43193, 43200, 43208, 43215, 43222, 43229, 43236, 43244, 43251, 43258, 43265, 43272, 43279, 43287, 43294, 43301, 43308, 43315, 43322, 43330, 43337, 43344, 43351, 43358, 43365, 43373, 43380, 43387, 43394, 43401, 43408, 43416, 43423, 43430, 43437, 43444, 43451, 43458, 43466, 43473, 43480, 43487, 43494, 43501, 43508, 43516, 43523, 43530, 43537, 43544, 43551, 43558, 43566, 43573, 43580, 43587, 43594, 43601, 43608, 43615, 43623, 43630, 43637, 43644, 43651, 43658, 43665, 43672, 43680, 43687, 43694, 43701, 43708, 43715, 43722, 43729, 43736, 43744, 43751, 43758, 43765, 43772, 43779, 43786, 43793, 43800, 43807, 43814, 43822, 43829, 43836, 43843, 43850, 43857, 43864, 43871, 43878, 43885, 43892, 43899, 43907, 43914, 43921, 43928, 43935, 43942, 43949, 43956, 43963, 43970, 43977, 43984, 43991, 43998, 44005, 44013, 44020, 44027, 44034, 44041, 44048, 44055, 44062, 44069, 44076, 44083, 44090, 44097, 44104, 44111, 44118, 44125, 44132, 44139, 44146, 44153, 44161, 44168, 44175, 44182, 44189, 44196, 44203, 44210, 44217, 44224, 44231, 44238, 44245, 44252, 44259, 44266, 44273, 44280, 44287, 44294, 44301, 44308, 44315, 44322, 44329, 44336, 44343, 44350, 44357, 44364, 44371, 44378, 44385, 44392, 44399, 44406, 44413, 44420, 44427, 44434, 44441, 44448, 44455, 44462, 44469, 44476, 44483, 44490, 44497, 44504, 44511, 44518, 44525, 44532, 44539, 44546, 44552, 44559, 44566, 44573, 44580, 44587, 44594, 44601, 44608, 44615, 44622, 44629, 44636, 44643, 44650, 44657, 44664, 44671, 44678, 44685, 44692, 44698, 44705, 44712, 44719, 44726, 44733, 44740, 44747, 44754, 44761, 44768, 44775, 44782, 44789, 44796, 44802, 44809, 44816, 44823, 44830, 44837, 44844, 44851, 44858, 44865, 44872, 44878, 44885, 44892, 44899, 44906, 44913, 44920, 44927, 44934, 44941, 44947, 44954, 44961, 44968, 44975, 44982, 44989, 44996, 45003, 45009, 45016, 45023, 45030, 45037, 45044, 45051, 45058, 45065, 45071, 45078, 45085, 45092, 45099, 45106, 45113, 45119, 45126, 45133, 45140, 45147, 45154, 45161, 45167, 45174, 45181, 45188, 45195, 45202, 45209, 45215, 45222, 45229, 45236, 45243, 45250, 45256, 45263, 45270, 45277, 45284, 45291, 45297, 45304, 45311, 45318, 45325, 45332, 45338, 45345, 45352, 45359, 45366, 45373, 45379, 45386, 45393, 45400, 45407, 45413, 45420, 45427, 45434, 45441, 45447, 45454, 45461, 45468, 45475, 45481, 45488, 45495, 45502, 45509, 45515, 45522, 45529, 45536, 45543, 45549, 45556, 45563, 45570, 45576, 45583, 45590, 45597, 45604, 45610, 45617, 45624, 45631, 45637, 45644, 45651, 45658, 45664, 45671, 45678, 45685, 45691, 45698, 45705, 45712, 45718, 45725, 45732, 45739, 45745, 45752, 45759, 45766, 45772, 45779, 45786, 45793, 45799, 45806, 45813, 45820, 45826, 45833, 45840, 45847, 45853, 45860, 45867, 45873, 45880, 45887, 45894, 45900, 45907, 45914, 45920, 45927, 45934, 45941, 45947, 45954, 45961, 45967, 45974, 45981, 45987, 45994, 46001, 46008, 46014, 46021, 46028, 46034, 46041, 46048, 46054, 46061, 46068, 46074, 46081, 46088, 46094, 46101, 46108, 46114, 46121, 46128, 46135, 46141, 46148, 46155, 46161, 46168, 46174, 46181, 46188, 46194, 46201, 46208, 46214, 46221, 46228, 46234, 46241, 46248, 46254, 46261, 46268, 46274, 46281, 46288, 46294, 46301, 46307, 46314, 46321, 46327, 46334, 46341, 46347, 46354, 46360, 46367, 46374, 46380, 46387, 46394, 46400, 46407, 46413, 46420, 46427, 46433, 46440, 46446, 46453, 46460, 46466, 46473, 46479, 46486, 46493, 46499, 46506, 46512, 46519, 46526, 46532, 46539, 46545, 46552, 46559, 46565, 46572, 46578, 46585, 46591, 46598, 46605, 46611, 46618, 46624, 46631, 46637, 46644, 46651, 46657, 46664, 46670, 46677, 46683, 46690, 46697, 46703, 46710, 46716, 46723, 46729, 46736, 46742, 46749, 46755, 46762, 46769, 46775, 46782, 46788, 46795, 46801, 46808, 46814, 46821, 46827, 46834, 46840, 46847, 46853, 46860, 46866, 46873, 46880, 46886, 46893, 46899, 46906, 46912, 46919, 46925, 46932, 46938, 46945, 46951, 46958, 46964, 46971, 46977, 46984, 46990, 46997, 47003, 47010, 47016, 47023, 47029, 47036, 47042, 47048, 47055, 47061, 47068, 47074, 47081, 47087, 47094, 47100, 47107, 47113, 47120, 47126, 47133, 47139, 47146, 47152, 47158, 47165, 47171, 47178, 47184, 47191, 47197, 47204, 47210, 47217, 47223, 47229, 47236, 47242, 47249, 47255, 47262, 47268, 47274, 47281, 47287, 47294, 47300, 47307, 47313, 47319, 47326, 47332, 47339, 47345, 47352, 47358, 47364, 47371, 47377, 47384, 47390, 47396, 47403, 47409, 47416, 47422, 47428, 47435, 47441, 47448, 47454, 47460, 47467, 47473, 47480, 47486, 47492, 47499, 47505, 47511, 47518, 47524, 47531, 47537, 47543, 47550, 47556, 47562, 47569, 47575, 47582, 47588, 47594, 47601, 47607, 47613, 47620, 47626, 47632, 47639, 47645, 47652, 47658, 47664, 47671, 47677, 47683, 47690, 47696, 47702, 47709, 47715, 47721, 47728, 47734, 47740, 47747, 47753, 47759, 47766, 47772, 47778, 47785, 47791, 47797, 47803, 47810, 47816, 47822, 47829, 47835, 47841, 47848, 47854, 47860, 47867, 47873, 47879, 47885, 47892, 47898, 47904, 47911, 47917, 47923, 47930, 47936, 47942, 47948, 47955, 47961, 47967, 47973, 47980, 47986, 47992, 47999, 48005, 48011, 48017, 48024, 48030, 48036, 48042, 48049, 48055, 48061, 48068, 48074, 48080, 48086, 48093, 48099, 48105, 48111, 48118, 48124, 48130, 48136, 48142, 48149, 48155, 48161, 48167, 48174, 48180, 48186, 48192, 48199, 48205, 48211, 48217, 48223, 48230, 48236, 48242, 48248, 48255, 48261, 48267, 48273, 48279, 48286, 48292, 48298, 48304, 48310, 48317, 48323, 48329, 48335, 48341, 48348, 48354, 48360, 48366, 48372, 48379, 48385, 48391, 48397, 48403, 48409, 48416, 48422, 48428, 48434, 48440, 48446, 48453, 48459, 48465, 48471, 48477, 48483, 48490, 48496, 48502, 48508, 48514, 48520, 48527, 48533, 48539, 48545, 48551, 48557, 48563, 48570, 48576, 48582, 48588, 48594, 48600, 48606, 48612, 48619, 48625, 48631, 48637, 48643, 48649, 48655, 48661, 48668, 48674, 48680, 48686, 48692, 48698, 48704, 48710, 48716, 48723, 48729, 48735, 48741, 48747, 48753, 48759, 48765, 48771, 48777, 48784, 48790, 48796, 48802, 48808, 48814, 48820, 48826, 48832, 48838, 48844, 48850, 48857, 48863, 48869, 48875, 48881, 48887, 48893, 48899, 48905, 48911, 48917, 48923, 48929, 48935, 48941, 48947, 48953, 48960, 48966, 48972, 48978, 48984, 48990, 48996, 49002, 49008, 49014, 49020, 49026, 49032, 49038, 49044, 49050, 49056, 49062, 49068, 49074, 49080, 49086, 49092, 49098, 49104, 49110, 49116, 49122, 49128, 49134, 49140, 49146, 49152, 49158, 49164, 49170, 49176, 49182, 49188, 49194, 49200, 49206, 49212, 49218, 49224, 49230, 49236, 49242, 49248, 49254, 49260, 49266, 49272, 49278, 49284, 49290, 49296, 49302, 49308, 49314, 49320, 49326, 49332, 49338, 49343, 49349, 49355, 49361, 49367, 49373, 49379, 49385, 49391, 49397, 49403, 49409, 49415, 49421, 49427, 49433, 49439, 49444, 49450, 49456, 49462, 49468, 49474, 49480, 49486, 49492, 49498, 49504, 49510, 49516, 49521, 49527, 49533, 49539, 49545, 49551, 49557, 49563, 49569, 49575, 49580, 49586, 49592, 49598, 49604, 49610, 49616, 49622, 49628, 49633, 49639, 49645, 49651, 49657, 49663, 49669, 49675, 49680, 49686, 49692, 49698, 49704, 49710, 49716, 49721, 49727, 49733, 49739, 49745, 49751, 49757, 49762, 49768, 49774, 49780, 49786, 49792, 49798, 49803, 49809, 49815, 49821, 49827, 49833, 49838, 49844, 49850, 49856, 49862, 49867, 49873, 49879, 49885, 49891, 49897, 49902, 49908, 49914, 49920, 49926, 49931, 49937, 49943, 49949, 49955, 49960, 49966, 49972, 49978, 49984, 49989, 49995, 50001, 50007, 50013, 50018, 50024, 50030, 50036, 50041, 50047, 50053, 50059, 50065, 50070, 50076, 50082, 50088, 50093, 50099, 50105, 50111, 50116, 50122, 50128, 50134, 50139, 50145, 50151, 50157, 50162, 50168, 50174, 50180, 50185, 50191, 50197, 50203, 50208, 50214, 50220, 50226, 50231, 50237, 50243, 50248, 50254, 50260, 50266, 50271, 50277, 50283, 50288, 50294, 50300, 50306, 50311, 50317, 50323, 50328, 50334, 50340, 50346, 50351, 50357, 50363, 50368, 50374, 50380, 50385, 50391, 50397, 50402, 50408, 50414, 50419, 50425, 50431, 50437, 50442, 50448, 50454, 50459, 50465, 50471, 50476, 50482, 50488, 50493, 50499, 50504, 50510, 50516, 50521, 50527, 50533, 50538, 50544, 50550, 50555, 50561, 50567, 50572, 50578, 50584, 50589, 50595, 50600, 50606, 50612, 50617, 50623, 50629, 50634, 50640, 50645, 50651, 50657, 50662, 50668, 50674, 50679, 50685, 50690, 50696, 50702, 50707, 50713, 50718, 50724, 50730, 50735, 50741, 50746, 50752, 50758, 50763, 50769, 50774, 50780, 50785, 50791, 50797, 50802, 50808, 50813, 50819, 50824, 50830, 50836, 50841, 50847, 50852, 50858, 50863, 50869, 50875, 50880, 50886, 50891, 50897, 50902, 50908, 50913, 50919, 50924, 50930, 50936, 50941, 50947, 50952, 50958, 50963, 50969, 50974, 50980, 50985, 50991, 50996, 51002, 51007, 51013, 51019, 51024, 51030, 51035, 51041, 51046, 51052, 51057, 51063, 51068, 51074, 51079, 51085, 51090, 51096, 51101, 51107, 51112, 51118, 51123, 51129, 51134, 51140, 51145, 51151, 51156, 51161, 51167, 51172, 51178, 51183, 51189, 51194, 51200, 51205, 51211, 51216, 51222, 51227, 51233, 51238, 51244, 51249, 51254, 51260, 51265, 51271, 51276, 51282, 51287, 51293, 51298, 51303, 51309, 51314, 51320, 51325, 51331, 51336, 51341, 51347, 51352, 51358, 51363, 51369, 51374, 51379, 51385, 51390, 51396, 51401, 51407, 51412, 51417, 51423, 51428, 51434, 51439, 51444, 51450, 51455, 51461, 51466, 51471, 51477, 51482, 51488, 51493, 51498, 51504, 51509, 51514, 51520, 51525, 51531, 51536, 51541, 51547, 51552, 51557, 51563, 51568, 51574, 51579, 51584, 51590, 51595, 51600, 51606, 51611, 51616, 51622, 51627, 51633, 51638, 51643, 51649, 51654, 51659, 51665, 51670, 51675, 51681, 51686, 51691, 51697, 51702, 51707, 51713, 51718, 51723, 51729, 51734, 51739, 51744, 51750, 51755, 51760, 51766, 51771, 51776, 51782, 51787, 51792, 51798, 51803, 51808, 51813, 51819, 51824, 51829, 51835, 51840, 51845, 51851, 51856, 51861, 51866, 51872, 51877, 51882, 51888, 51893, 51898, 51903, 51909, 51914, 51919, 51924, 51930, 51935, 51940, 51945, 51951, 51956, 51961, 51966, 51972, 51977, 51982, 51987, 51993, 51998, 52003, 52008, 52014, 52019, 52024, 52029, 52035, 52040, 52045, 52050, 52056, 52061, 52066, 52071, 52076, 52082, 52087, 52092, 52097, 52103, 52108, 52113, 52118, 52123, 52129, 52134, 52139, 52144, 52149, 52155, 52160, 52165, 52170, 52175, 52181, 52186, 52191, 52196, 52201, 52207, 52212, 52217, 52222, 52227, 52232, 52238, 52243, 52248, 52253, 52258, 52264, 52269, 52274, 52279, 52284, 52289, 52294, 52300, 52305, 52310, 52315, 52320, 52325, 52331, 52336, 52341, 52346, 52351, 52356, 52361, 52367, 52372, 52377, 52382, 52387, 52392, 52397, 52403, 52408, 52413, 52418, 52423, 52428, 52433, 52438, 52443, 52449, 52454, 52459, 52464, 52469, 52474, 52479, 52484, 52489, 52495, 52500, 52505, 52510, 52515, 52520, 52525, 52530, 52535, 52540, 52545, 52551, 52556, 52561, 52566, 52571, 52576, 52581, 52586, 52591, 52596, 52601, 52606, 52611, 52617, 52622, 52627, 52632, 52637, 52642, 52647, 52652, 52657, 52662, 52667, 52672, 52677, 52682, 52687, 52692, 52697, 52702, 52707, 52713, 52718, 52723, 52728, 52733, 52738, 52743, 52748, 52753, 52758, 52763, 52768, 52773, 52778, 52783, 52788, 52793, 52798, 52803, 52808, 52813, 52818, 52823, 52828, 52833, 52838, 52843, 52848, 52853, 52858, 52863, 52868, 52873, 52878, 52883, 52888, 52893, 52898, 52903, 52908, 52913, 52918, 52923, 52928, 52933, 52938, 52943, 52948, 52953, 52957, 52962, 52967, 52972, 52977, 52982, 52987, 52992, 52997, 53002, 53007, 53012, 53017, 53022, 53027, 53032, 53037, 53042, 53047, 53052, 53056, 53061, 53066, 53071, 53076, 53081, 53086, 53091, 53096, 53101, 53106, 53111, 53116, 53120, 53125, 53130, 53135, 53140, 53145, 53150, 53155, 53160, 53165, 53170, 53174, 53179, 53184, 53189, 53194, 53199, 53204, 53209, 53214, 53218, 53223, 53228, 53233, 53238, 53243, 53248, 53253, 53257, 53262, 53267, 53272, 53277, 53282, 53287, 53292, 53296, 53301, 53306, 53311, 53316, 53321, 53326, 53330, 53335, 53340, 53345, 53350, 53355, 53359, 53364, 53369, 53374, 53379, 53384, 53388, 53393, 53398, 53403, 53408, 53413, 53417, 53422, 53427, 53432, 53437, 53442, 53446, 53451, 53456, 53461, 53466, 53470, 53475, 53480, 53485, 53490, 53494, 53499, 53504, 53509, 53514, 53518, 53523, 53528, 53533, 53538, 53542, 53547, 53552, 53557, 53561, 53566, 53571, 53576, 53581, 53585, 53590, 53595, 53600, 53604, 53609, 53614, 53619, 53623, 53628, 53633, 53638, 53642, 53647, 53652, 53657, 53661, 53666, 53671, 53676, 53680, 53685, 53690, 53695, 53699, 53704, 53709, 53714, 53718, 53723, 53728, 53733, 53737, 53742, 53747, 53751, 53756, 53761, 53766, 53770, 53775, 53780, 53784, 53789, 53794, 53799, 53803, 53808, 53813, 53817, 53822, 53827, 53831, 53836, 53841, 53846, 53850, 53855, 53860, 53864, 53869, 53874, 53878, 53883, 53888, 53892, 53897, 53902, 53906, 53911, 53916, 53920, 53925, 53930, 53934, 53939, 53944, 53948, 53953, 53958, 53962, 53967, 53972, 53976, 53981, 53986, 53990, 53995, 53999, 54004, 54009, 54013, 54018, 54023, 54027, 54032, 54037, 54041, 54046, 54050, 54055, 54060, 54064, 54069, 54074, 54078, 54083, 54087, 54092, 54097, 54101, 54106, 54110, 54115, 54120, 54124, 54129, 54133, 54138, 54143, 54147, 54152, 54156, 54161, 54166, 54170, 54175, 54179, 54184, 54189, 54193, 54198, 54202, 54207, 54211, 54216, 54221, 54225, 54230, 54234, 54239, 54243, 54248, 54253, 54257, 54262, 54266, 54271, 54275, 54280, 54284, 54289, 54294, 54298, 54303, 54307, 54312, 54316, 54321, 54325, 54330, 54334, 54339, 54343, 54348, 54353, 54357, 54362, 54366, 54371, 54375, 54380, 54384, 54389, 54393, 54398, 54402, 54407, 54411, 54416, 54420, 54425, 54429, 54434, 54438, 54443, 54447, 54452, 54456, 54461, 54465, 54470, 54474, 54479, 54483, 54488, 54492, 54497, 54501, 54506, 54510, 54515, 54519, 54524, 54528, 54533, 54537, 54541, 54546, 54550, 54555, 54559, 54564, 54568, 54573, 54577, 54582, 54586, 54591, 54595, 54599, 54604, 54608, 54613, 54617, 54622, 54626, 54631, 54635, 54639, 54644, 54648, 54653, 54657, 54662, 54666, 54670, 54675, 54679, 54684, 54688, 54693, 54697, 54701, 54706, 54710, 54715, 54719, 54723, 54728, 54732, 54737, 54741, 54745, 54750, 54754, 54759, 54763, 54767, 54772, 54776, 54781, 54785, 54789, 54794, 54798, 54803, 54807, 54811, 54816, 54820, 54824, 54829, 54833, 54838, 54842, 54846, 54851, 54855, 54859, 54864, 54868, 54872, 54877, 54881, 54886, 54890, 54894, 54899, 54903, 54907, 54912, 54916, 54920, 54925, 54929, 54933, 54938, 54942, 54946, 54951, 54955, 54959, 54964, 54968, 54972, 54977, 54981, 54985, 54990, 54994, 54998, 55003, 55007, 55011, 55016, 55020, 55024, 55028, 55033, 55037, 55041, 55046, 55050, 55054, 55059, 55063, 55067, 55072, 55076, 55080, 55084, 55089, 55093, 55097, 55102, 55106, 55110, 55114, 55119, 55123, 55127, 55131, 55136, 55140, 55144, 55149, 55153, 55157, 55161, 55166, 55170, 55174, 55178, 55183, 55187, 55191, 55195, 55200, 55204, 55208, 55212, 55217, 55221, 55225, 55229, 55234, 55238, 55242, 55246, 55251, 55255, 55259, 55263, 55268, 55272, 55276, 55280, 55284, 55289, 55293, 55297, 55301, 55306, 55310, 55314, 55318, 55322, 55327, 55331, 55335, 55339, 55343, 55348, 55352, 55356, 55360, 55364, 55369, 55373, 55377, 55381, 55385, 55390, 55394, 55398, 55402, 55406, 55410, 55415, 55419, 55423, 55427, 55431, 55436, 55440, 55444, 55448, 55452, 55456, 55461, 55465, 55469, 55473, 55477, 55481, 55485, 55490, 55494, 55498, 55502, 55506, 55510, 55515, 55519, 55523, 55527, 55531, 55535, 55539, 55544, 55548, 55552, 55556, 55560, 55564, 55568, 55572, 55577, 55581, 55585, 55589, 55593, 55597, 55601, 55605, 55609, 55614, 55618, 55622, 55626, 55630, 55634, 55638, 55642, 55646, 55651, 55655, 55659, 55663, 55667, 55671, 55675, 55679, 55683, 55687, 55691, 55696, 55700, 55704, 55708, 55712, 55716, 55720, 55724, 55728, 55732, 55736, 55740, 55744, 55749, 55753, 55757, 55761, 55765, 55769, 55773, 55777, 55781, 55785, 55789, 55793, 55797, 55801, 55805, 55809, 55813, 55817, 55821, 55826, 55830, 55834, 55838, 55842, 55846, 55850, 55854, 55858, 55862, 55866, 55870, 55874, 55878, 55882, 55886, 55890, 55894, 55898, 55902, 55906, 55910, 55914, 55918, 55922, 55926, 55930, 55934, 55938, 55942, 55946, 55950, 55954, 55958, 55962, 55966, 55970, 55974, 55978, 55982, 55986, 55990, 55994, 55998, 56002, 56006, 56010, 56014, 56018, 56022, 56026, 56030, 56034, 56038, 56042, 56046, 56050, 56053, 56057, 56061, 56065, 56069, 56073, 56077, 56081, 56085, 56089, 56093, 56097, 56101, 56105, 56109, 56113, 56117, 56121, 56125, 56128, 56132, 56136, 56140, 56144, 56148, 56152, 56156, 56160, 56164, 56168, 56172, 56176, 56179, 56183, 56187, 56191, 56195, 56199, 56203, 56207, 56211, 56215, 56219, 56222, 56226, 56230, 56234, 56238, 56242, 56246, 56250, 56254, 56258, 56261, 56265, 56269, 56273, 56277, 56281, 56285, 56289, 56292, 56296, 56300, 56304, 56308, 56312, 56316, 56320, 56323, 56327, 56331, 56335, 56339, 56343, 56347, 56350, 56354, 56358, 56362, 56366, 56370, 56374, 56377, 56381, 56385, 56389, 56393, 56397, 56401, 56404, 56408, 56412, 56416, 56420, 56424, 56427, 56431, 56435, 56439, 56443, 56446, 56450, 56454, 56458, 56462, 56466, 56469, 56473, 56477, 56481, 56485, 56488, 56492, 56496, 56500, 56504, 56507, 56511, 56515, 56519, 56523, 56526, 56530, 56534, 56538, 56542, 56545, 56549, 56553, 56557, 56561, 56564, 56568, 56572, 56576, 56579, 56583, 56587, 56591, 56595, 56598, 56602, 56606, 56610, 56613, 56617, 56621, 56625, 56628, 56632, 56636, 56640, 56643, 56647, 56651, 56655, 56658, 56662, 56666, 56670, 56673, 56677, 56681, 56685, 56688, 56692, 56696, 56700, 56703, 56707, 56711, 56715, 56718, 56722, 56726, 56729, 56733, 56737, 56741, 56744, 56748, 56752, 56755, 56759, 56763, 56767, 56770, 56774, 56778, 56781, 56785, 56789, 56793, 56796, 56800, 56804, 56807, 56811, 56815, 56818, 56822, 56826, 56829, 56833, 56837, 56840, 56844, 56848, 56852, 56855, 56859, 56863, 56866, 56870, 56874, 56877, 56881, 56885, 56888, 56892, 56896, 56899, 56903, 56907, 56910, 56914, 56918, 56921, 56925, 56928, 56932, 56936, 56939, 56943, 56947, 56950, 56954, 56958, 56961, 56965, 56969, 56972, 56976, 56979, 56983, 56987, 56990, 56994, 56998, 57001, 57005, 57008, 57012, 57016, 57019, 57023, 57027, 57030, 57034, 57037, 57041, 57045, 57048, 57052, 57055, 57059, 57063, 57066, 57070, 57073, 57077, 57081, 57084, 57088, 57091, 57095, 57099, 57102, 57106, 57109, 57113, 57117, 57120, 57124, 57127, 57131, 57134, 57138, 57142, 57145, 57149, 57152, 57156, 57159, 57163, 57167, 57170, 57174, 57177, 57181, 57184, 57188, 57192, 57195, 57199, 57202, 57206, 57209, 57213, 57216, 57220, 57223, 57227, 57231, 57234, 57238, 57241, 57245, 57248, 57252, 57255, 57259, 57262, 57266, 57269, 57273, 57276, 57280, 57284, 57287, 57291, 57294, 57298, 57301, 57305, 57308, 57312, 57315, 57319, 57322, 57326, 57329, 57333, 57336, 57340, 57343, 57347, 57350, 57354, 57357, 57361, 57364, 57368, 57371, 57375, 57378, 57382, 57385, 57389, 57392, 57396, 57399, 57403, 57406, 57409, 57413, 57416, 57420, 57423, 57427, 57430, 57434, 57437, 57441, 57444, 57448, 57451, 57455, 57458, 57461, 57465, 57468, 57472, 57475, 57479, 57482, 57486, 57489, 57493, 57496, 57499, 57503, 57506, 57510, 57513, 57517, 57520, 57524, 57527, 57530, 57534, 57537, 57541, 57544, 57548, 57551, 57554, 57558, 57561, 57565, 57568, 57571, 57575, 57578, 57582, 57585, 57589, 57592, 57595, 57599, 57602, 57606, 57609, 57612, 57616, 57619, 57623, 57626, 57629, 57633, 57636, 57640, 57643, 57646, 57650, 57653, 57656, 57660, 57663, 57667, 57670, 57673, 57677, 57680, 57684, 57687, 57690, 57694, 57697, 57700, 57704, 57707, 57710, 57714, 57717, 57721, 57724, 57727, 57731, 57734, 57737, 57741, 57744, 57747, 57751, 57754, 57757, 57761, 57764, 57767, 57771, 57774, 57778, 57781, 57784, 57788, 57791, 57794, 57798, 57801, 57804, 57808, 57811, 57814, 57818, 57821, 57824, 57827, 57831, 57834, 57837, 57841, 57844, 57847, 57851, 57854, 57857, 57861, 57864, 57867, 57871, 57874, 57877, 57880, 57884, 57887, 57890, 57894, 57897, 57900, 57904, 57907, 57910, 57913, 57917, 57920, 57923, 57927, 57930, 57933, 57936, 57940, 57943, 57946, 57950, 57953, 57956, 57959, 57963, 57966, 57969, 57972, 57976, 57979, 57982, 57985, 57989, 57992, 57995, 57999, 58002, 58005, 58008, 58012, 58015, 58018, 58021, 58025, 58028, 58031, 58034, 58038, 58041, 58044, 58047, 58050, 58054, 58057, 58060, 58063, 58067, 58070, 58073, 58076, 58080, 58083, 58086, 58089, 58092, 58096, 58099, 58102, 58105, 58109, 58112, 58115, 58118, 58121, 58125, 58128, 58131, 58134, 58137, 58141, 58144, 58147, 58150, 58153, 58157, 58160, 58163, 58166, 58169, 58173, 58176, 58179, 58182, 58185, 58189, 58192, 58195, 58198, 58201, 58204, 58208, 58211, 58214, 58217, 58220, 58224, 58227, 58230, 58233, 58236, 58239, 58243, 58246, 58249, 58252, 58255, 58258, 58261, 58265, 58268, 58271, 58274, 58277, 58280, 58284, 58287, 58290, 58293, 58296, 58299, 58302, 58306, 58309, 58312, 58315, 58318, 58321, 58324, 58328, 58331, 58334, 58337, 58340, 58343, 58346, 58349, 58353, 58356, 58359, 58362, 58365, 58368, 58371, 58374, 58378, 58381, 58384, 58387, 58390, 58393, 58396, 58399, 58402, 58405, 58409, 58412, 58415, 58418, 58421, 58424, 58427, 58430, 58433, 58436, 58440, 58443, 58446, 58449, 58452, 58455, 58458, 58461, 58464, 58467, 58470, 58473, 58477, 58480, 58483, 58486, 58489, 58492, 58495, 58498, 58501, 58504, 58507, 58510, 58513, 58516, 58519, 58523, 58526, 58529, 58532, 58535, 58538, 58541, 58544, 58547, 58550, 58553, 58556, 58559, 58562, 58565, 58568, 58571, 58574, 58577, 58580, 58583, 58587, 58590, 58593, 58596, 58599, 58602, 58605, 58608, 58611, 58614, 58617, 58620, 58623, 58626, 58629, 58632, 58635, 58638, 58641, 58644, 58647, 58650, 58653, 58656, 58659, 58662, 58665, 58668, 58671, 58674, 58677, 58680, 58683, 58686, 58689, 58692, 58695, 58698, 58701, 58704, 58707, 58710, 58713, 58716, 58719, 58722, 58725, 58728, 58731, 58734, 58737, 58740, 58743, 58746, 58749, 58752, 58755, 58758, 58760, 58763, 58766, 58769, 58772, 58775, 58778, 58781, 58784, 58787, 58790, 58793, 58796, 58799, 58802, 58805, 58808, 58811, 58814, 58817, 58820, 58823, 58825, 58828, 58831, 58834, 58837, 58840, 58843, 58846, 58849, 58852, 58855, 58858, 58861, 58864, 58867, 58869, 58872, 58875, 58878, 58881, 58884, 58887, 58890, 58893, 58896, 58899, 58902, 58904, 58907, 58910, 58913, 58916, 58919, 58922, 58925, 58928, 58931, 58934, 58936, 58939, 58942, 58945, 58948, 58951, 58954, 58957, 58960, 58962, 58965, 58968, 58971, 58974, 58977, 58980, 58983, 58986, 58988, 58991, 58994, 58997, 59000, 59003, 59006, 59009, 59011, 59014, 59017, 59020, 59023, 59026, 59029, 59031, 59034, 59037, 59040, 59043, 59046, 59049, 59051, 59054, 59057, 59060, 59063, 59066, 59069, 59071, 59074, 59077, 59080, 59083, 59086, 59088, 59091, 59094, 59097, 59100, 59103, 59105, 59108, 59111, 59114, 59117, 59120, 59122, 59125, 59128, 59131, 59134, 59137, 59139, 59142, 59145, 59148, 59151, 59153, 59156, 59159, 59162, 59165, 59167, 59170, 59173, 59176, 59179, 59181, 59184, 59187, 59190, 59193, 59195, 59198, 59201, 59204, 59207, 59209, 59212, 59215, 59218, 59221, 59223, 59226, 59229, 59232, 59235, 59237, 59240, 59243, 59246, 59248, 59251, 59254, 59257, 59260, 59262, 59265, 59268, 59271, 59273, 59276, 59279, 59282, 59284, 59287, 59290, 59293, 59295, 59298, 59301, 59304, 59306, 59309, 59312, 59315, 59317, 59320, 59323, 59326, 59328, 59331, 59334, 59337, 59339, 59342, 59345, 59348, 59350, 59353, 59356, 59359, 59361, 59364, 59367, 59369, 59372, 59375, 59378, 59380, 59383, 59386, 59389, 59391, 59394, 59397, 59399, 59402, 59405, 59408, 59410, 59413, 59416, 59418, 59421, 59424, 59427, 59429, 59432, 59435, 59437, 59440, 59443, 59445, 59448, 59451, 59454, 59456, 59459, 59462, 59464, 59467, 59470, 59472, 59475, 59478, 59480, 59483, 59486, 59488, 59491, 59494, 59497, 59499, 59502, 59505, 59507, 59510, 59513, 59515, 59518, 59521, 59523, 59526, 59529, 59531, 59534, 59537, 59539, 59542, 59545, 59547, 59550, 59552, 59555, 59558, 59560, 59563, 59566, 59568, 59571, 59574, 59576, 59579, 59582, 59584, 59587, 59590, 59592, 59595, 59597, 59600, 59603, 59605, 59608, 59611, 59613, 59616, 59619, 59621, 59624, 59626, 59629, 59632, 59634, 59637, 59640, 59642, 59645, 59647, 59650, 59653, 59655, 59658, 59660, 59663, 59666, 59668, 59671, 59674, 59676, 59679, 59681, 59684, 59687, 59689, 59692, 59694, 59697, 59700, 59702, 59705, 59707, 59710, 59712, 59715, 59718, 59720, 59723, 59725, 59728, 59731, 59733, 59736, 59738, 59741, 59743, 59746, 59749, 59751, 59754, 59756, 59759, 59762, 59764, 59767, 59769, 59772, 59774, 59777, 59779, 59782, 59785, 59787, 59790, 59792, 59795, 59797, 59800, 59803, 59805, 59808, 59810, 59813, 59815, 59818, 59820, 59823, 59825, 59828, 59831, 59833, 59836, 59838, 59841, 59843, 59846, 59848, 59851, 59853, 59856, 59858, 59861, 59864, 59866, 59869, 59871, 59874, 59876, 59879, 59881, 59884, 59886, 59889, 59891, 59894, 59896, 59899, 59901, 59904, 59906, 59909, 59911, 59914, 59916, 59919, 59921, 59924, 59926, 59929, 59931, 59934, 59936, 59939, 59941, 59944, 59946, 59949, 59951, 59954, 59956, 59959, 59961, 59964, 59966, 59969, 59971, 59974, 59976, 59979, 59981, 59984, 59986, 59989, 59991, 59994, 59996, 59999, 60001, 60004, 60006, 60009, 60011, 60014, 60016, 60018, 60021, 60023, 60026, 60028, 60031, 60033, 60036, 60038, 60041, 60043, 60046, 60048, 60050, 60053, 60055, 60058, 60060, 60063, 60065, 60068, 60070, 60072, 60075, 60077, 60080, 60082, 60085, 60087, 60090, 60092, 60094, 60097, 60099, 60102, 60104, 60107, 60109, 60111, 60114, 60116, 60119, 60121, 60124, 60126, 60128, 60131, 60133, 60136, 60138, 60141, 60143, 60145, 60148, 60150, 60153, 60155, 60157, 60160, 60162, 60165, 60167, 60170, 60172, 60174, 60177, 60179, 60182, 60184, 60186, 60189, 60191, 60194, 60196, 60198, 60201, 60203, 60205, 60208, 60210, 60213, 60215, 60217, 60220, 60222, 60225, 60227, 60229, 60232, 60234, 60236, 60239, 60241, 60244, 60246, 60248, 60251, 60253, 60255, 60258, 60260, 60263, 60265, 60267, 60270, 60272, 60274, 60277, 60279, 60282, 60284, 60286, 60289, 60291, 60293, 60296, 60298, 60300, 60303, 60305, 60307, 60310, 60312, 60314, 60317, 60319, 60321, 60324, 60326, 60329, 60331, 60333, 60336, 60338, 60340, 60343, 60345, 60347, 60350, 60352, 60354, 60357, 60359, 60361, 60364, 60366, 60368, 60370, 60373, 60375, 60377, 60380, 60382, 60384, 60387, 60389, 60391, 60394, 60396, 60398, 60401, 60403, 60405, 60408, 60410, 60412, 60414, 60417, 60419, 60421, 60424, 60426, 60428, 60431, 60433, 60435, 60437, 60440, 60442, 60444, 60447, 60449, 60451, 60454, 60456, 60458, 60460, 60463, 60465, 60467, 60470, 60472, 60474, 60476, 60479, 60481, 60483, 60485, 60488, 60490, 60492, 60495, 60497, 60499, 60501, 60504, 60506, 60508, 60510, 60513, 60515, 60517, 60520, 60522, 60524, 60526, 60529, 60531, 60533, 60535, 60538, 60540, 60542, 60544, 60547, 60549, 60551, 60553, 60556, 60558, 60560, 60562, 60565, 60567, 60569, 60571, 60574, 60576, 60578, 60580, 60582, 60585, 60587, 60589, 60591, 60594, 60596, 60598, 60600, 60603, 60605, 60607, 60609, 60611, 60614, 60616, 60618, 60620, 60623, 60625, 60627, 60629, 60631, 60634, 60636, 60638, 60640, 60643, 60645, 60647, 60649, 60651, 60654, 60656, 60658, 60660, 60662, 60665, 60667, 60669, 60671, 60673, 60676, 60678, 60680, 60682, 60684, 60687, 60689, 60691, 60693, 60695, 60697, 60700, 60702, 60704, 60706, 60708, 60711, 60713, 60715, 60717, 60719, 60722, 60724, 60726, 60728, 60730, 60732, 60735, 60737, 60739, 60741, 60743, 60745, 60748, 60750, 60752, 60754, 60756, 60758, 60761, 60763, 60765, 60767, 60769, 60771, 60774, 60776, 60778, 60780, 60782, 60784, 60786, 60789, 60791, 60793, 60795, 60797, 60799, 60801, 60804, 60806, 60808, 60810, 60812, 60814, 60816, 60819, 60821, 60823, 60825, 60827, 60829, 60831, 60834, 60836, 60838, 60840, 60842, 60844, 60846, 60848, 60851, 60853, 60855, 60857, 60859, 60861, 60863, 60865, 60868, 60870, 60872, 60874, 60876, 60878, 60880, 60882, 60884, 60887, 60889, 60891, 60893, 60895, 60897, 60899, 60901, 60903, 60906, 60908, 60910, 60912, 60914, 60916, 60918, 60920, 60922, 60924, 60926, 60929, 60931, 60933, 60935, 60937, 60939, 60941, 60943, 60945, 60947, 60949, 60952, 60954, 60956, 60958, 60960, 60962, 60964, 60966, 60968, 60970, 60972, 60974, 60976, 60979, 60981, 60983, 60985, 60987, 60989, 60991, 60993, 60995, 60997, 60999, 61001, 61003, 61005, 61007, 61009, 61012, 61014, 61016, 61018, 61020, 61022, 61024, 61026, 61028, 61030, 61032, 61034, 61036, 61038, 61040, 61042, 61044, 61046, 61048, 61050, 61052, 61055, 61057, 61059, 61061, 61063, 61065, 61067, 61069, 61071, 61073, 61075, 61077, 61079, 61081, 61083, 61085, 61087, 61089, 61091, 61093, 61095, 61097, 61099, 61101, 61103, 61105, 61107, 61109, 61111, 61113, 61115, 61117, 61119, 61121, 61123, 61125, 61127, 61129, 61131, 61133, 61135, 61137, 61139, 61141, 61143, 61145, 61147, 61149, 61151, 61153, 61155, 61157, 61159, 61161, 61163, 61165, 61167, 61169, 61171, 61173, 61175, 61177, 61179, 61181, 61183, 61185, 61187, 61189, 61191, 61193, 61195, 61197, 61199, 61201, 61203, 61205, 61207, 61209, 61211, 61213, 61215, 61217, 61219, 61221, 61223, 61225, 61227, 61229, 61231, 61233, 61235, 61237, 61238, 61240, 61242, 61244, 61246, 61248, 61250, 61252, 61254, 61256, 61258, 61260, 61262, 61264, 61266, 61268, 61270, 61272, 61274, 61276, 61278, 61279, 61281, 61283, 61285, 61287, 61289, 61291, 61293, 61295, 61297, 61299, 61301, 61303, 61305, 61307, 61309, 61310, 61312, 61314, 61316, 61318, 61320, 61322, 61324, 61326, 61328, 61330, 61332, 61334, 61335, 61337, 61339, 61341, 61343, 61345, 61347, 61349, 61351, 61353, 61355, 61357, 61358, 61360, 61362, 61364, 61366, 61368, 61370, 61372, 61374, 61376, 61378, 61379, 61381, 61383, 61385, 61387, 61389, 61391, 61393, 61395, 61396, 61398, 61400, 61402, 61404, 61406, 61408, 61410, 61412, 61414, 61415, 61417, 61419, 61421, 61423, 61425, 61427, 61429, 61430, 61432, 61434, 61436, 61438, 61440, 61442, 61444, 61445, 61447, 61449, 61451, 61453, 61455, 61457, 61459, 61460, 61462, 61464, 61466, 61468, 61470, 61472, 61473, 61475, 61477, 61479, 61481, 61483, 61485, 61486, 61488, 61490, 61492, 61494, 61496, 61498, 61499, 61501, 61503, 61505, 61507, 61509, 61511, 61512, 61514, 61516, 61518, 61520, 61522, 61523, 61525, 61527, 61529, 61531, 61533, 61534, 61536, 61538, 61540, 61542, 61544, 61545, 61547, 61549, 61551, 61553, 61555, 61556, 61558, 61560, 61562, 61564, 61566, 61567, 61569, 61571, 61573, 61575, 61576, 61578, 61580, 61582, 61584, 61585, 61587, 61589, 61591, 61593, 61595, 61596, 61598, 61600, 61602, 61604, 61605, 61607, 61609, 61611, 61613, 61614, 61616, 61618, 61620, 61622, 61623, 61625, 61627, 61629, 61631, 61632, 61634, 61636, 61638, 61640, 61641, 61643, 61645, 61647, 61648, 61650, 61652, 61654, 61656, 61657, 61659, 61661, 61663, 61665, 61666, 61668, 61670, 61672, 61673, 61675, 61677, 61679, 61680, 61682, 61684, 61686, 61688, 61689, 61691, 61693, 61695, 61696, 61698, 61700, 61702, 61703, 61705, 61707, 61709, 61710, 61712, 61714, 61716, 61718, 61719, 61721, 61723, 61725, 61726, 61728, 61730, 61732, 61733, 61735, 61737, 61739, 61740, 61742, 61744, 61746, 61747, 61749, 61751, 61752, 61754, 61756, 61758, 61759, 61761, 61763, 61765, 61766, 61768, 61770, 61772, 61773, 61775, 61777, 61779, 61780, 61782, 61784, 61785, 61787, 61789, 61791, 61792, 61794, 61796, 61797, 61799, 61801, 61803, 61804, 61806, 61808, 61810, 61811, 61813, 61815, 61816, 61818, 61820, 61822, 61823, 61825, 61827, 61828, 61830, 61832, 61833, 61835, 61837, 61839, 61840, 61842, 61844, 61845, 61847, 61849, 61850, 61852, 61854, 61856, 61857, 61859, 61861, 61862, 61864, 61866, 61867, 61869, 61871, 61873, 61874, 61876, 61878, 61879, 61881, 61883, 61884, 61886, 61888, 61889, 61891, 61893, 61894, 61896, 61898, 61899, 61901, 61903, 61904, 61906, 61908, 61909, 61911, 61913, 61915, 61916, 61918, 61920, 61921, 61923, 61925, 61926, 61928, 61930, 61931, 61933, 61934, 61936, 61938, 61939, 61941, 61943, 61944, 61946, 61948, 61949, 61951, 61953, 61954, 61956, 61958, 61959, 61961, 61963, 61964, 61966, 61968, 61969, 61971, 61973, 61974, 61976, 61977, 61979, 61981, 61982, 61984, 61986, 61987, 61989, 61991, 61992, 61994, 61995, 61997, 61999, 62000, 62002, 62004, 62005, 62007, 62009, 62010, 62012, 62013, 62015, 62017, 62018, 62020, 62022, 62023, 62025, 62026, 62028, 62030, 62031, 62033, 62035, 62036, 62038, 62039, 62041, 62043, 62044, 62046, 62047, 62049, 62051, 62052, 62054, 62056, 62057, 62059, 62060, 62062, 62064, 62065, 62067, 62068, 62070, 62072, 62073, 62075, 62076, 62078, 62080, 62081, 62083, 62084, 62086, 62088, 62089, 62091, 62092, 62094, 62096, 62097, 62099, 62100, 62102, 62103, 62105, 62107, 62108, 62110, 62111, 62113, 62115, 62116, 62118, 62119, 62121, 62122, 62124, 62126, 62127, 62129, 62130, 62132, 62134, 62135, 62137, 62138, 62140, 62141, 62143, 62145, 62146, 62148, 62149, 62151, 62152, 62154, 62156, 62157, 62159, 62160, 62162, 62163, 62165, 62166, 62168, 62170, 62171, 62173, 62174, 62176, 62177, 62179, 62180, 62182, 62184, 62185, 62187, 62188, 62190, 62191, 62193, 62194, 62196, 62198, 62199, 62201, 62202, 62204, 62205, 62207, 62208, 62210, 62211, 62213, 62215, 62216, 62218, 62219, 62221, 62222, 62224, 62225, 62227, 62228, 62230, 62231, 62233, 62234, 62236, 62238, 62239, 62241, 62242, 62244, 62245, 62247, 62248, 62250, 62251, 62253, 62254, 62256, 62257, 62259, 62260, 62262, 62263, 62265, 62266, 62268, 62270, 62271, 62273, 62274, 62276, 62277, 62279, 62280, 62282, 62283, 62285, 62286, 62288, 62289, 62291, 62292, 62294, 62295, 62297, 62298, 62300, 62301, 62303, 62304, 62306, 62307, 62309, 62310, 62312, 62313, 62315, 62316, 62318, 62319, 62321, 62322, 62324, 62325, 62327, 62328, 62330, 62331, 62333, 62334, 62336, 62337, 62339, 62340, 62341, 62343, 62344, 62346, 62347, 62349, 62350, 62352, 62353, 62355, 62356, 62358, 62359, 62361, 62362, 62364, 62365, 62367, 62368, 62370, 62371, 62372, 62374, 62375, 62377, 62378, 62380, 62381, 62383, 62384, 62386, 62387, 62389, 62390, 62392, 62393, 62394, 62396, 62397, 62399, 62400, 62402, 62403, 62405, 62406, 62408, 62409, 62411, 62412, 62413, 62415, 62416, 62418, 62419, 62421, 62422, 62424, 62425, 62426, 62428, 62429, 62431, 62432, 62434, 62435, 62437, 62438, 62439, 62441, 62442, 62444, 62445, 62447, 62448, 62450, 62451, 62452, 62454, 62455, 62457, 62458, 62460, 62461, 62462, 62464, 62465, 62467, 62468, 62470, 62471, 62472, 62474, 62475, 62477, 62478, 62480, 62481, 62482, 62484, 62485, 62487, 62488, 62489, 62491, 62492, 62494, 62495, 62497, 62498, 62499, 62501, 62502, 62504, 62505, 62506, 62508, 62509, 62511, 62512, 62513, 62515, 62516, 62518, 62519, 62521, 62522, 62523, 62525, 62526, 62528, 62529, 62530, 62532, 62533, 62535, 62536, 62537, 62539, 62540, 62542, 62543, 62544, 62546, 62547, 62548, 62550, 62551, 62553, 62554, 62555, 62557, 62558, 62560, 62561, 62562, 62564, 62565, 62567, 62568, 62569, 62571, 62572, 62573, 62575, 62576, 62578, 62579, 62580, 62582, 62583, 62584, 62586, 62587, 62589, 62590, 62591, 62593, 62594, 62595, 62597, 62598, 62600, 62601, 62602, 62604, 62605, 62606, 62608, 62609, 62611, 62612, 62613, 62615, 62616, 62617, 62619, 62620, 62621, 62623, 62624, 62626, 62627, 62628, 62630, 62631, 62632, 62634, 62635, 62636, 62638, 62639, 62640, 62642, 62643, 62644, 62646, 62647, 62648, 62650, 62651, 62653, 62654, 62655, 62657, 62658, 62659, 62661, 62662, 62663, 62665, 62666, 62667, 62669, 62670, 62671, 62673, 62674, 62675, 62677, 62678, 62679, 62681, 62682, 62683, 62685, 62686, 62687, 62689, 62690, 62691, 62693, 62694, 62695, 62697, 62698, 62699, 62701, 62702, 62703, 62705, 62706, 62707, 62709, 62710, 62711, 62713, 62714, 62715, 62716, 62718, 62719, 62720, 62722, 62723, 62724, 62726, 62727, 62728, 62730, 62731, 62732, 62734, 62735, 62736, 62737, 62739, 62740, 62741, 62743, 62744, 62745, 62747, 62748, 62749, 62751, 62752, 62753, 62754, 62756, 62757, 62758, 62760, 62761, 62762, 62764, 62765, 62766, 62767, 62769, 62770, 62771, 62773, 62774, 62775, 62776, 62778, 62779, 62780, 62782, 62783, 62784, 62785, 62787, 62788, 62789, 62791, 62792, 62793, 62794, 62796, 62797, 62798, 62800, 62801, 62802, 62803, 62805, 62806, 62807, 62809, 62810, 62811, 62812, 62814, 62815, 62816, 62817, 62819, 62820, 62821, 62823, 62824, 62825, 62826, 62828, 62829, 62830, 62831, 62833, 62834, 62835, 62836, 62838, 62839, 62840, 62842, 62843, 62844, 62845, 62847, 62848, 62849, 62850, 62852, 62853, 62854, 62855, 62857, 62858, 62859, 62860, 62862, 62863, 62864, 62865, 62867, 62868, 62869, 62870, 62872, 62873, 62874, 62875, 62877, 62878, 62879, 62880, 62882, 62883, 62884, 62885, 62887, 62888, 62889, 62890, 62892, 62893, 62894, 62895, 62896, 62898, 62899, 62900, 62901, 62903, 62904, 62905, 62906, 62908, 62909, 62910, 62911, 62913, 62914, 62915, 62916, 62917, 62919, 62920, 62921, 62922, 62924, 62925, 62926, 62927, 62928, 62930, 62931, 62932, 62933, 62935, 62936, 62937, 62938, 62939, 62941, 62942, 62943, 62944, 62946, 62947, 62948, 62949, 62950, 62952, 62953, 62954, 62955, 62956, 62958, 62959, 62960, 62961, 62962, 62964, 62965, 62966, 62967, 62969, 62970, 62971, 62972, 62973, 62975, 62976, 62977, 62978, 62979, 62981, 62982, 62983, 62984, 62985, 62987, 62988, 62989, 62990, 62991, 62992, 62994, 62995, 62996, 62997, 62998, 63000, 63001, 63002, 63003, 63004, 63006, 63007, 63008, 63009, 63010, 63012, 63013, 63014, 63015, 63016, 63017, 63019, 63020, 63021, 63022, 63023, 63025, 63026, 63027, 63028, 63029, 63030, 63032, 63033, 63034, 63035, 63036, 63037, 63039, 63040, 63041, 63042, 63043, 63045, 63046, 63047, 63048, 63049, 63050, 63052, 63053, 63054, 63055, 63056, 63057, 63059, 63060, 63061, 63062, 63063, 63064, 63065, 63067, 63068, 63069, 63070, 63071, 63072, 63074, 63075, 63076, 63077, 63078, 63079, 63081, 63082, 63083, 63084, 63085, 63086, 63087, 63089, 63090, 63091, 63092, 63093, 63094, 63095, 63097, 63098, 63099, 63100, 63101, 63102, 63104, 63105, 63106, 63107, 63108, 63109, 63110, 63111, 63113, 63114, 63115, 63116, 63117, 63118, 63119, 63121, 63122, 63123, 63124, 63125, 63126, 63127, 63129, 63130, 63131, 63132, 63133, 63134, 63135, 63136, 63138, 63139, 63140, 63141, 63142, 63143, 63144, 63145, 63147, 63148, 63149, 63150, 63151, 63152, 63153, 63154, 63156, 63157, 63158, 63159, 63160, 63161, 63162, 63163, 63165, 63166, 63167, 63168, 63169, 63170, 63171, 63172, 63173, 63175, 63176, 63177, 63178, 63179, 63180, 63181, 63182, 63183, 63185, 63186, 63187, 63188, 63189, 63190, 63191, 63192, 63193, 63194, 63196, 63197, 63198, 63199, 63200, 63201, 63202, 63203, 63204, 63205, 63207, 63208, 63209, 63210, 63211, 63212, 63213, 63214, 63215, 63216, 63218, 63219, 63220, 63221, 63222, 63223, 63224, 63225, 63226, 63227, 63228, 63229, 63231, 63232, 63233, 63234, 63235, 63236, 63237, 63238, 63239, 63240, 63241, 63242, 63244, 63245, 63246, 63247, 63248, 63249, 63250, 63251, 63252, 63253, 63254, 63255, 63257, 63258, 63259, 63260, 63261, 63262, 63263, 63264, 63265, 63266, 63267, 63268, 63269, 63270, 63271, 63273, 63274, 63275, 63276, 63277, 63278, 63279, 63280, 63281, 63282, 63283, 63284, 63285, 63286, 63287, 63289, 63290, 63291, 63292, 63293, 63294, 63295, 63296, 63297, 63298, 63299, 63300, 63301, 63302, 63303, 63304, 63305, 63306, 63308, 63309, 63310, 63311, 63312, 63313, 63314, 63315, 63316, 63317, 63318, 63319, 63320, 63321, 63322, 63323, 63324, 63325, 63326, 63327, 63328, 63329, 63331, 63332, 63333, 63334, 63335, 63336, 63337, 63338, 63339, 63340, 63341, 63342, 63343, 63344, 63345, 63346, 63347, 63348, 63349, 63350, 63351, 63352, 63353, 63354, 63355, 63356, 63357, 63358, 63359, 63360, 63362, 63363, 63364, 63365, 63366, 63367, 63368, 63369, 63370, 63371, 63372, 63373, 63374, 63375, 63376, 63377, 63378, 63379, 63380, 63381, 63382, 63383, 63384, 63385, 63386, 63387, 63388, 63389, 63390, 63391, 63392, 63393, 63394, 63395, 63396, 63397, 63398, 63399, 63400, 63401, 63402, 63403, 63404, 63405, 63406, 63407, 63408, 63409, 63410, 63411, 63412, 63413, 63414, 63415, 63416, 63417, 63418, 63419, 63420, 63421, 63422, 63423, 63424, 63425, 63426, 63427, 63428, 63429, 63430, 63431, 63432, 63433, 63434, 63435, 63436, 63437, 63438, 63439, 63440, 63441, 63442, 63443, 63444, 63445, 63446, 63447, 63448, 63449, 63450, 63451, 63452, 63453, 63454, 63455, 63456, 63457, 63458, 63459, 63460, 63461, 63462, 63463, 63464, 63465, 63466, 63467, 63468, 63469, 63470, 63471, 63472, 63473, 63474, 63475, 63476, 63477, 63478, 63478, 63479, 63480, 63481, 63482, 63483, 63484, 63485, 63486, 63487, 63488, 63489, 63490, 63491, 63492, 63493, 63494, 63495, 63496, 63497, 63498, 63499, 63500, 63501, 63502, 63503, 63504, 63505, 63506, 63507, 63507, 63508, 63509, 63510, 63511, 63512, 63513, 63514, 63515, 63516, 63517, 63518, 63519, 63520, 63521, 63522, 63523, 63524, 63525, 63526, 63527, 63528, 63528, 63529, 63530, 63531, 63532, 63533, 63534, 63535, 63536, 63537, 63538, 63539, 63540, 63541, 63542, 63543, 63544, 63545, 63546, 63546, 63547, 63548, 63549, 63550, 63551, 63552, 63553, 63554, 63555, 63556, 63557, 63558, 63559, 63560, 63561, 63561, 63562, 63563, 63564, 63565, 63566, 63567, 63568, 63569, 63570, 63571, 63572, 63573, 63574, 63575, 63575, 63576, 63577, 63578, 63579, 63580, 63581, 63582, 63583, 63584, 63585, 63586, 63587, 63587, 63588, 63589, 63590, 63591, 63592, 63593, 63594, 63595, 63596, 63597, 63598, 63599, 63599, 63600, 63601, 63602, 63603, 63604, 63605, 63606, 63607, 63608, 63609, 63610, 63610, 63611, 63612, 63613, 63614, 63615, 63616, 63617, 63618, 63619, 63620, 63620, 63621, 63622, 63623, 63624, 63625, 63626, 63627, 63628, 63629, 63630, 63630, 63631, 63632, 63633, 63634, 63635, 63636, 63637, 63638, 63639, 63639, 63640, 63641, 63642, 63643, 63644, 63645, 63646, 63647, 63648, 63648, 63649, 63650, 63651, 63652, 63653, 63654, 63655, 63656, 63656, 63657, 63658, 63659, 63660, 63661, 63662, 63663, 63664, 63664, 63665, 63666, 63667, 63668, 63669, 63670, 63671, 63672, 63672, 63673, 63674, 63675, 63676, 63677, 63678, 63679, 63679, 63680, 63681, 63682, 63683, 63684, 63685, 63686, 63687, 63687, 63688, 63689, 63690, 63691, 63692, 63693, 63694, 63694, 63695, 63696, 63697, 63698, 63699, 63700, 63700, 63701, 63702, 63703, 63704, 63705, 63706, 63707, 63707, 63708, 63709, 63710, 63711, 63712, 63713, 63714, 63714, 63715, 63716, 63717, 63718, 63719, 63720, 63720, 63721, 63722, 63723, 63724, 63725, 63726, 63726, 63727, 63728, 63729, 63730, 63731, 63732, 63732, 63733, 63734, 63735, 63736, 63737, 63738, 63738, 63739, 63740, 63741, 63742, 63743, 63744, 63744, 63745, 63746, 63747, 63748, 63749, 63750, 63750, 63751, 63752, 63753, 63754, 63755, 63755, 63756, 63757, 63758, 63759, 63760, 63761, 63761, 63762, 63763, 63764, 63765, 63766, 63766, 63767, 63768, 63769, 63770, 63771, 63771, 63772, 63773, 63774, 63775, 63776, 63776, 63777, 63778, 63779, 63780, 63781, 63781, 63782, 63783, 63784, 63785, 63786, 63786, 63787, 63788, 63789, 63790, 63791, 63791, 63792, 63793, 63794, 63795, 63796, 63796, 63797, 63798, 63799, 63800, 63801, 63801, 63802, 63803, 63804, 63805, 63805, 63806, 63807, 63808, 63809, 63810, 63810, 63811, 63812, 63813, 63814, 63815, 63815, 63816, 63817, 63818, 63819, 63819, 63820, 63821, 63822, 63823, 63823, 63824, 63825, 63826, 63827, 63828, 63828, 63829, 63830, 63831, 63832, 63832, 63833, 63834, 63835, 63836, 63836, 63837, 63838, 63839, 63840, 63841, 63841, 63842, 63843, 63844, 63845, 63845, 63846, 63847, 63848, 63849, 63849, 63850, 63851, 63852, 63853, 63853, 63854, 63855, 63856, 63857, 63857, 63858, 63859, 63860, 63861, 63861, 63862, 63863, 63864, 63865, 63865, 63866, 63867, 63868, 63869, 63869, 63870, 63871, 63872, 63872, 63873, 63874, 63875, 63876, 63876, 63877, 63878, 63879, 63880, 63880, 63881, 63882, 63883, 63884, 63884, 63885, 63886, 63887, 63887, 63888, 63889, 63890, 63891, 63891, 63892, 63893, 63894, 63894, 63895, 63896, 63897, 63898, 63898, 63899, 63900, 63901, 63902, 63902, 63903, 63904, 63905, 63905, 63906, 63907, 63908, 63909, 63909, 63910, 63911, 63912, 63912, 63913, 63914, 63915, 63915, 63916, 63917, 63918, 63919, 63919, 63920, 63921, 63922, 63922, 63923, 63924, 63925, 63925, 63926, 63927, 63928, 63929, 63929, 63930, 63931, 63932, 63932, 63933, 63934, 63935, 63935, 63936, 63937, 63938, 63938, 63939, 63940, 63941, 63941, 63942, 63943, 63944, 63945, 63945, 63946, 63947, 63948, 63948, 63949, 63950, 63951, 63951, 63952, 63953, 63954, 63954, 63955, 63956, 63957, 63957, 63958, 63959, 63960, 63960, 63961, 63962, 63963, 63963, 63964, 63965, 63966, 63966, 63967, 63968, 63969, 63969, 63970, 63971, 63972, 63972, 63973, 63974, 63975, 63975, 63976, 63977, 63978, 63978, 63979, 63980, 63981, 63981, 63982, 63983, 63983, 63984, 63985, 63986, 63986, 63987, 63988, 63989, 63989, 63990, 63991, 63992, 63992, 63993, 63994, 63995, 63995, 63996, 63997, 63997, 63998, 63999, 64000, 64000, 64001, 64002, 64003, 64003, 64004, 64005, 64006, 64006, 64007, 64008, 64008, 64009, 64010, 64011, 64011, 64012, 64013, 64014, 64014, 64015, 64016, 64016, 64017, 64018, 64019, 64019, 64020, 64021, 64022, 64022, 64023, 64024, 64024, 64025, 64026, 64027, 64027, 64028, 64029, 64029, 64030, 64031, 64032, 64032, 64033, 64034, 64034, 64035, 64036, 64037, 64037, 64038, 64039, 64039, 64040, 64041, 64042, 64042, 64043, 64044, 64044, 64045, 64046, 64047, 64047, 64048, 64049, 64049, 64050, 64051, 64052, 64052, 64053, 64054, 64054, 64055, 64056, 64057, 64057, 64058, 64059, 64059, 64060, 64061, 64061, 64062, 64063, 64064, 64064, 64065, 64066, 64066, 64067, 64068, 64068, 64069, 64070, 64071, 64071, 64072, 64073, 64073, 64074, 64075, 64075, 64076, 64077, 64078, 64078, 64079, 64080, 64080, 64081, 64082, 64082, 64083, 64084, 64084, 64085, 64086, 64087, 64087, 64088, 64089, 64089, 64090, 64091, 64091, 64092, 64093, 64093, 64094, 64095, 64096, 64096, 64097, 64098, 64098, 64099, 64100, 64100, 64101, 64102, 64102, 64103, 64104, 64104, 64105, 64106, 64107, 64107, 64108, 64109, 64109, 64110, 64111, 64111, 64112, 64113, 64113, 64114, 64115, 64115, 64116, 64117, 64117, 64118, 64119, 64119, 64120, 64121, 64121, 64122, 64123, 64123, 64124, 64125, 64125, 64126, 64127, 64128, 64128, 64129, 64130, 64130, 64131, 64132, 64132, 64133, 64134, 64134, 64135, 64136, 64136, 64137, 64138, 64138, 64139, 64140, 64140, 64141, 64142, 64142, 64143, 64144, 64144, 64145, 64146, 64146, 64147, 64148, 64148, 64149, 64150, 64150, 64151, 64152, 64152, 64153, 64154, 64154, 64155, 64156, 64156, 64157, 64157, 64158, 64159, 64159, 64160, 64161, 64161, 64162, 64163, 64163, 64164, 64165, 64165, 64166, 64167, 64167, 64168, 64169, 64169, 64170, 64171, 64171, 64172, 64173, 64173, 64174, 64175, 64175, 64176, 64176, 64177, 64178, 64178, 64179, 64180, 64180, 64181, 64182, 64182, 64183, 64184, 64184, 64185, 64186, 64186, 64187, 64187, 64188, 64189, 64189, 64190, 64191, 64191, 64192, 64193, 64193, 64194, 64195, 64195, 64196, 64196, 64197, 64198, 64198, 64199, 64200, 64200, 64201, 64202, 64202, 64203, 64203, 64204, 64205, 64205, 64206, 64207, 64207, 64208, 64209, 64209, 64210, 64210, 64211, 64212, 64212, 64213, 64214, 64214, 64215, 64216, 64216, 64217, 64217, 64218, 64219, 64219, 64220, 64221, 64221, 64222, 64222, 64223, 64224, 64224, 64225, 64226, 64226, 64227, 64228, 64228, 64229, 64229, 64230, 64231, 64231, 64232, 64233, 64233, 64234, 64234, 64235, 64236, 64236, 64237, 64237, 64238, 64239, 64239, 64240, 64241, 64241, 64242, 64242, 64243, 64244, 64244, 64245, 64246, 64246, 64247, 64247, 64248, 64249, 64249, 64250, 64250, 64251, 64252, 64252, 64253, 64254, 64254, 64255, 64255, 64256, 64257, 64257, 64258, 64258, 64259, 64260, 64260, 64261, 64262, 64262, 64263, 64263, 64264, 64265, 64265, 64266, 64266, 64267, 64268, 64268, 64269, 64269, 64270, 64271, 64271, 64272, 64272, 64273, 64274, 64274, 64275, 64275, 64276, 64277, 64277, 64278, 64278, 64279, 64280, 64280, 64281, 64281, 64282, 64283, 64283, 64284, 64284, 64285, 64286, 64286, 64287, 64287, 64288, 64289, 64289, 64290, 64290, 64291, 64292, 64292, 64293, 64293, 64294, 64295, 64295, 64296, 64296, 64297, 64298, 64298, 64299, 64299, 64300, 64301, 64301, 64302, 64302, 64303, 64304, 64304, 64305, 64305, 64306, 64306, 64307, 64308, 64308, 64309, 64309, 64310, 64311, 64311, 64312, 64312, 64313, 64314, 64314, 64315, 64315, 64316, 64316, 64317, 64318, 64318, 64319, 64319, 64320, 64321, 64321, 64322, 64322, 64323, 64323, 64324, 64325, 64325, 64326, 64326, 64327, 64328, 64328, 64329, 64329, 64330, 64330, 64331, 64332, 64332, 64333, 64333, 64334, 64334, 64335, 64336, 64336, 64337, 64337, 64338, 64338, 64339, 64340, 64340, 64341, 64341, 64342, 64342, 64343, 64344, 64344, 64345, 64345, 64346, 64346, 64347, 64348, 64348, 64349, 64349, 64350, 64350, 64351, 64352, 64352, 64353, 64353, 64354, 64354, 64355, 64356, 64356, 64357, 64357, 64358, 64358, 64359, 64360, 64360, 64361, 64361, 64362, 64362, 64363, 64363, 64364, 64365, 64365, 64366, 64366, 64367, 64367, 64368, 64369, 64369, 64370, 64370, 64371, 64371, 64372, 64372, 64373, 64374, 64374, 64375, 64375, 64376, 64376, 64377, 64377, 64378, 64379, 64379, 64380, 64380, 64381, 64381, 64382, 64382, 64383, 64384, 64384, 64385, 64385, 64386, 64386, 64387, 64387, 64388, 64388, 64389, 64390, 64390, 64391, 64391, 64392, 64392, 64393, 64393, 64394, 64395, 64395, 64396, 64396, 64397, 64397, 64398, 64398, 64399, 64399, 64400, 64401, 64401, 64402, 64402, 64403, 64403, 64404, 64404, 64405, 64405, 64406, 64407, 64407, 64408, 64408, 64409, 64409, 64410, 64410, 64411, 64411, 64412, 64412, 64413, 64414, 64414, 64415, 64415, 64416, 64416, 64417, 64417, 64418, 64418, 64419, 64419, 64420, 64421, 64421, 64422, 64422, 64423, 64423, 64424, 64424, 64425, 64425, 64426, 64426, 64427, 64427, 64428, 64429, 64429, 64430, 64430, 64431, 64431, 64432, 64432, 64433, 64433, 64434, 64434, 64435, 64435, 64436, 64436, 64437, 64438, 64438, 64439, 64439, 64440, 64440, 64441, 64441, 64442, 64442, 64443, 64443, 64444, 64444, 64445, 64445, 64446, 64446, 64447, 64448, 64448, 64449, 64449, 64450, 64450, 64451, 64451, 64452, 64452, 64453, 64453, 64454, 64454, 64455, 64455, 64456, 64456, 64457, 64457, 64458, 64458, 64459, 64459, 64460, 64460, 64461, 64462, 64462, 64463, 64463, 64464, 64464, 64465, 64465, 64466, 64466, 64467, 64467, 64468, 64468, 64469, 64469, 64470, 64470, 64471, 64471, 64472, 64472, 64473, 64473, 64474, 64474, 64475, 64475, 64476, 64476, 64477, 64477, 64478, 64478, 64479, 64479, 64480, 64480, 64481, 64481, 64482, 64482, 64483, 64483, 64484, 64485, 64485, 64486, 64486, 64487, 64487, 64488, 64488, 64489, 64489, 64490, 64490, 64491, 64491, 64492, 64492, 64493, 64493, 64494, 64494, 64495, 64495, 64496, 64496, 64497, 64497, 64498, 64498, 64499, 64499, 64500, 64500, 64501, 64501, 64502, 64502, 64503, 64503, 64504, 64504, 64505, 64505, 64506, 64506, 64507, 64507, 64507, 64508, 64508, 64509, 64509, 64510, 64510, 64511, 64511, 64512, 64512, 64513, 64513, 64514, 64514, 64515, 64515, 64516, 64516, 64517, 64517, 64518, 64518, 64519, 64519, 64520, 64520, 64521, 64521, 64522, 64522, 64523, 64523, 64524, 64524, 64525, 64525, 64526, 64526, 64527, 64527, 64528, 64528, 64529, 64529, 64530, 64530, 64530, 64531, 64531, 64532, 64532, 64533, 64533, 64534, 64534, 64535, 64535, 64536, 64536, 64537, 64537, 64538, 64538, 64539, 64539, 64540, 64540, 64541, 64541, 64542, 64542, 64542, 64543, 64543, 64544, 64544, 64545, 64545, 64546, 64546, 64547, 64547, 64548, 64548, 64549, 64549, 64550, 64550, 64551, 64551, 64552, 64552, 64552, 64553, 64553, 64554, 64554, 64555, 64555, 64556, 64556, 64557, 64557, 64558, 64558, 64559, 64559, 64560, 64560, 64560, 64561, 64561, 64562, 64562, 64563, 64563, 64564, 64564, 64565, 64565, 64566, 64566, 64567, 64567, 64567, 64568, 64568, 64569, 64569, 64570, 64570, 64571, 64571, 64572, 64572, 64573, 64573, 64574, 64574, 64574, 64575, 64575, 64576, 64576, 64577, 64577, 64578, 64578, 64579, 64579, 64580, 64580, 64580, 64581, 64581, 64582, 64582, 64583, 64583, 64584, 64584, 64585, 64585, 64585, 64586, 64586, 64587, 64587, 64588, 64588, 64589, 64589, 64590, 64590, 64591, 64591, 64591, 64592, 64592, 64593, 64593, 64594, 64594, 64595, 64595, 64596, 64596, 64596, 64597, 64597, 64598, 64598, 64599, 64599, 64600, 64600, 64600, 64601, 64601, 64602, 64602, 64603, 64603, 64604, 64604, 64605, 64605, 64605, 64606, 64606, 64607, 64607, 64608, 64608, 64609, 64609, 64609, 64610, 64610, 64611, 64611, 64612, 64612, 64613, 64613, 64613, 64614, 64614, 64615, 64615, 64616, 64616, 64617, 64617, 64617, 64618, 64618, 64619, 64619, 64620, 64620, 64621, 64621, 64621, 64622, 64622, 64623, 64623, 64624, 64624, 64624, 64625, 64625, 64626, 64626, 64627, 64627, 64628, 64628, 64628, 64629, 64629, 64630, 64630, 64631, 64631, 64631, 64632, 64632, 64633, 64633, 64634, 64634, 64635, 64635, 64635, 64636, 64636, 64637, 64637, 64638, 64638, 64638, 64639, 64639, 64640, 64640, 64641, 64641, 64641, 64642, 64642, 64643, 64643, 64644, 64644, 64644, 64645, 64645, 64646, 64646, 64647, 64647, 64647, 64648, 64648, 64649, 64649, 64650, 64650, 64650, 64651, 64651, 64652, 64652, 64653, 64653, 64653, 64654, 64654, 64655, 64655, 64656, 64656, 64656, 64657, 64657, 64658, 64658, 64659, 64659, 64659, 64660, 64660, 64661, 64661, 64661, 64662, 64662, 64663, 64663, 64664, 64664, 64664, 64665, 64665, 64666, 64666, 64667, 64667, 64667, 64668, 64668, 64669, 64669, 64669, 64670, 64670, 64671, 64671, 64672, 64672, 64672, 64673, 64673, 64674, 64674, 64674, 64675, 64675, 64676, 64676, 64676, 64677, 64677, 64678, 64678, 64679, 64679, 64679, 64680, 64680, 64681, 64681, 64681, 64682, 64682, 64683, 64683, 64684, 64684, 64684, 64685, 64685, 64686, 64686, 64686, 64687, 64687, 64688, 64688, 64688, 64689, 64689, 64690, 64690, 64690, 64691, 64691, 64692, 64692, 64693, 64693, 64693, 64694, 64694, 64695, 64695, 64695, 64696, 64696, 64697, 64697, 64697, 64698, 64698, 64699, 64699, 64699, 64700, 64700, 64701, 64701, 64701, 64702, 64702, 64703, 64703, 64703, 64704, 64704, 64705, 64705, 64705, 64706, 64706, 64707, 64707, 64707, 64708, 64708, 64709, 64709, 64709, 64710, 64710, 64711, 64711, 64711, 64712, 64712, 64713, 64713, 64713, 64714, 64714, 64715, 64715, 64715, 64716, 64716, 64717, 64717, 64717, 64718, 64718, 64719, 64719, 64719, 64720, 64720, 64720, 64721, 64721, 64722, 64722, 64722, 64723, 64723, 64724, 64724, 64724, 64725, 64725, 64726, 64726, 64726, 64727, 64727, 64728, 64728, 64728, 64729, 64729, 64729, 64730, 64730, 64731, 64731, 64731, 64732, 64732, 64733, 64733, 64733, 64734, 64734, 64735, 64735, 64735, 64736, 64736, 64736, 64737, 64737, 64738, 64738, 64738, 64739, 64739, 64740, 64740, 64740, 64741, 64741, 64741, 64742, 64742, 64743, 64743, 64743, 64744, 64744, 64745, 64745, 64745, 64746, 64746, 64746, 64747, 64747, 64748, 64748, 64748, 64749, 64749, 64749, 64750, 64750, 64751, 64751, 64751, 64752, 64752, 64752, 64753, 64753, 64754, 64754, 64754, 64755, 64755, 64756, 64756, 64756, 64757, 64757, 64757, 64758, 64758, 64759, 64759, 64759, 64760, 64760, 64760, 64761, 64761, 64762, 64762, 64762, 64763, 64763, 64763, 64764, 64764, 64764, 64765, 64765, 64766, 64766, 64766, 64767, 64767, 64767, 64768, 64768, 64769, 64769, 64769, 64770, 64770, 64770, 64771, 64771, 64772, 64772, 64772, 64773, 64773, 64773, 64774, 64774, 64774, 64775, 64775, 64776, 64776, 64776, 64777, 64777, 64777, 64778, 64778, 64779, 64779, 64779, 64780, 64780, 64780, 64781, 64781, 64781, 64782, 64782, 64783, 64783, 64783, 64784, 64784, 64784, 64785, 64785, 64785, 64786, 64786, 64787, 64787, 64787, 64788, 64788, 64788, 64789, 64789, 64789, 64790, 64790, 64790, 64791, 64791, 64792, 64792, 64792, 64793, 64793, 64793, 64794, 64794, 64794, 64795, 64795, 64796, 64796, 64796, 64797, 64797, 64797, 64798, 64798, 64798, 64799, 64799, 64799, 64800, 64800, 64800, 64801, 64801, 64802, 64802, 64802, 64803, 64803, 64803, 64804, 64804, 64804, 64805, 64805, 64805, 64806, 64806, 64807, 64807, 64807, 64808, 64808, 64808, 64809, 64809, 64809, 64810, 64810, 64810, 64811, 64811, 64811, 64812, 64812, 64812, 64813, 64813, 64814, 64814, 64814, 64815, 64815, 64815, 64816, 64816, 64816, 64817, 64817, 64817, 64818, 64818, 64818, 64819, 64819, 64819, 64820, 64820, 64820, 64821, 64821, 64822, 64822, 64822, 64823, 64823, 64823, 64824, 64824, 64824, 64825, 64825, 64825, 64826, 64826, 64826, 64827, 64827, 64827, 64828, 64828, 64828, 64829, 64829, 64829, 64830, 64830, 64830, 64831, 64831, 64831, 64832, 64832, 64832, 64833, 64833, 64833, 64834, 64834, 64834, 64835, 64835, 64836, 64836, 64836, 64837, 64837, 64837, 64838, 64838, 64838, 64839, 64839, 64839, 64840, 64840, 64840, 64841, 64841, 64841, 64842, 64842, 64842, 64843, 64843, 64843, 64844, 64844, 64844, 64845, 64845, 64845, 64846, 64846, 64846, 64847, 64847, 64847, 64848, 64848, 64848, 64849, 64849, 64849, 64850, 64850, 64850, 64851, 64851, 64851, 64852, 64852, 64852, 64853, 64853, 64853, 64854, 64854, 64854, 64855, 64855, 64855, 64856, 64856, 64856, 64857, 64857, 64857, 64857, 64858, 64858, 64858, 64859, 64859, 64859, 64860, 64860, 64860, 64861, 64861, 64861, 64862, 64862, 64862, 64863, 64863, 64863, 64864, 64864, 64864, 64865, 64865, 64865, 64866, 64866, 64866, 64867, 64867, 64867, 64868, 64868, 64868, 64869, 64869, 64869, 64870, 64870, 64870, 64870, 64871, 64871, 64871, 64872, 64872, 64872, 64873, 64873, 64873, 64874, 64874, 64874, 64875, 64875, 64875, 64876, 64876, 64876, 64877, 64877, 64877, 64878, 64878, 64878, 64878, 64879, 64879, 64879, 64880, 64880, 64880, 64881, 64881, 64881, 64882, 64882, 64882, 64883, 64883, 64883, 64884, 64884, 64884, 64884, 64885, 64885, 64885, 64886, 64886, 64886, 64887, 64887, 64887, 64888, 64888, 64888, 64889, 64889, 64889, 64890, 64890, 64890, 64890, 64891, 64891, 64891, 64892, 64892, 64892, 64893, 64893, 64893, 64894, 64894, 64894, 64894, 64895, 64895, 64895, 64896, 64896, 64896, 64897, 64897, 64897, 64898, 64898, 64898, 64899, 64899, 64899, 64899, 64900, 64900, 64900, 64901, 64901, 64901, 64902, 64902, 64902, 64903, 64903, 64903, 64903, 64904, 64904, 64904, 64905, 64905, 64905, 64906, 64906, 64906, 64906, 64907, 64907, 64907, 64908, 64908, 64908, 64909, 64909, 64909, 64910, 64910, 64910, 64910, 64911, 64911, 64911, 64912, 64912, 64912, 64913, 64913, 64913, 64913, 64914, 64914, 64914, 64915, 64915, 64915, 64916, 64916, 64916, 64916, 64917, 64917, 64917, 64918, 64918, 64918, 64919, 64919, 64919, 64919, 64920, 64920, 64920, 64921, 64921, 64921, 64922, 64922, 64922, 64922, 64923, 64923, 64923, 64924, 64924, 64924, 64924, 64925, 64925, 64925, 64926, 64926, 64926, 64927, 64927, 64927, 64927, 64928, 64928, 64928, 64929, 64929, 64929, 64929, 64930, 64930, 64930, 64931, 64931, 64931, 64932, 64932, 64932, 64932, 64933, 64933, 64933, 64934, 64934, 64934, 64934, 64935, 64935, 64935, 64936, 64936, 64936, 64936, 64937, 64937, 64937, 64938, 64938, 64938, 64939, 64939, 64939, 64939, 64940, 64940, 64940, 64941, 64941, 64941, 64941, 64942, 64942, 64942, 64943, 64943, 64943, 64943, 64944, 64944, 64944, 64945, 64945, 64945, 64945, 64946, 64946, 64946, 64947, 64947, 64947, 64947, 64948, 64948, 64948, 64949, 64949, 64949, 64949, 64950, 64950, 64950, 64951, 64951, 64951, 64951, 64952, 64952, 64952, 64953, 64953, 64953, 64953, 64954, 64954, 64954, 64954, 64955, 64955, 64955, 64956, 64956, 64956, 64956, 64957, 64957, 64957, 64958, 64958, 64958, 64958, 64959, 64959, 64959, 64960, 64960, 64960, 64960, 64961, 64961, 64961, 64961, 64962, 64962, 64962, 64963, 64963, 64963, 64963, 64964, 64964, 64964, 64965, 64965, 64965, 64965, 64966, 64966, 64966, 64966, 64967, 64967, 64967, 64968, 64968, 64968, 64968, 64969, 64969, 64969, 64969, 64970, 64970, 64970, 64971, 64971, 64971, 64971, 64972, 64972, 64972, 64973, 64973, 64973, 64973, 64974, 64974, 64974, 64974, 64975, 64975, 64975, 64975, 64976, 64976, 64976, 64977, 64977, 64977, 64977, 64978, 64978, 64978, 64978, 64979, 64979, 64979, 64980, 64980, 64980, 64980, 64981, 64981, 64981, 64981, 64982, 64982, 64982, 64983, 64983, 64983, 64983, 64984, 64984, 64984, 64984, 64985, 64985, 64985, 64985, 64986, 64986, 64986, 64987, 64987, 64987, 64987, 64988, 64988, 64988, 64988, 64989, 64989, 64989, 64989, 64990, 64990, 64990, 64990, 64991, 64991, 64991, 64992, 64992, 64992, 64992, 64993, 64993, 64993, 64993, 64994, 64994, 64994, 64994, 64995, 64995, 64995, 64995, 64996, 64996, 64996, 64997, 64997, 64997, 64997, 64998, 64998, 64998, 64998, 64999, 64999, 64999, 64999, 65000, 65000, 65000, 65000, 65001, 65001, 65001, 65001, 65002, 65002, 65002, 65003, 65003, 65003, 65003, 65004, 65004, 65004, 65004, 65005, 65005, 65005, 65005, 65006, 65006, 65006, 65006, 65007, 65007, 65007, 65007, 65008, 65008, 65008, 65008, 65009, 65009, 65009, 65009, 65010, 65010, 65010, 65010, 65011, 65011, 65011, 65011, 65012, 65012, 65012, 65012, 65013, 65013, 65013, 65014, 65014, 65014, 65014, 65015, 65015, 65015, 65015, 65016, 65016, 65016, 65016, 65017, 65017, 65017, 65017, 65018, 65018, 65018, 65018, 65019, 65019, 65019, 65019, 65020, 65020, 65020, 65020, 65021, 65021, 65021, 65021, 65022, 65022, 65022, 65022, 65023, 65023, 65023, 65023, 65024, 65024, 65024, 65024, 65025, 65025, 65025, 65025, 65026, 65026, 65026, 65026, 65027, 65027, 65027, 65027, 65027, 65028, 65028, 65028, 65028, 65029, 65029, 65029, 65029, 65030, 65030, 65030, 65030, 65031, 65031, 65031, 65031, 65032, 65032, 65032, 65032, 65033, 65033, 65033, 65033, 65034, 65034, 65034, 65034, 65035, 65035, 65035, 65035, 65036, 65036, 65036, 65036, 65037, 65037, 65037, 65037, 65037, 65038, 65038, 65038, 65038, 65039, 65039, 65039, 65039, 65040, 65040, 65040, 65040, 65041, 65041, 65041, 65041, 65042, 65042, 65042, 65042, 65043, 65043, 65043, 65043, 65043, 65044, 65044, 65044, 65044, 65045, 65045, 65045, 65045, 65046, 65046, 65046, 65046, 65047, 65047, 65047, 65047, 65048, 65048, 65048, 65048, 65048, 65049, 65049, 65049, 65049, 65050, 65050, 65050, 65050, 65051, 65051, 65051, 65051, 65052, 65052, 65052, 65052, 65052, 65053, 65053, 65053, 65053, 65054, 65054, 65054, 65054, 65055, 65055, 65055, 65055, 65056, 65056, 65056, 65056, 65056, 65057, 65057, 65057, 65057, 65058, 65058, 65058, 65058, 65059, 65059, 65059, 65059, 65059, 65060, 65060, 65060, 65060, 65061, 65061, 65061, 65061, 65062, 65062, 65062, 65062, 65062, 65063, 65063, 65063, 65063, 65064, 65064, 65064, 65064, 65065, 65065, 65065, 65065, 65065, 65066, 65066, 65066, 65066, 65067, 65067, 65067, 65067, 65067, 65068, 65068, 65068, 65068, 65069, 65069, 65069, 65069, 65070, 65070, 65070, 65070, 65070, 65071, 65071, 65071, 65071, 65072, 65072, 65072, 65072, 65072, 65073, 65073, 65073, 65073, 65074, 65074, 65074, 65074, 65074, 65075, 65075, 65075, 65075, 65076, 65076, 65076, 65076, 65076, 65077, 65077, 65077, 65077, 65078, 65078, 65078, 65078, 65078, 65079, 65079, 65079, 65079, 65080, 65080, 65080, 65080, 65080, 65081, 65081, 65081, 65081, 65082, 65082, 65082, 65082, 65082, 65083, 65083, 65083, 65083, 65084, 65084, 65084, 65084, 65084, 65085, 65085, 65085, 65085, 65086, 65086, 65086, 65086, 65086, 65087, 65087, 65087, 65087, 65087, 65088, 65088, 65088, 65088, 65089, 65089, 65089, 65089, 65089, 65090, 65090, 65090, 65090, 65091, 65091, 65091, 65091, 65091, 65092, 65092, 65092, 65092, 65092, 65093, 65093, 65093, 65093, 65094, 65094, 65094, 65094, 65094, 65095, 65095, 65095, 65095, 65095, 65096, 65096, 65096, 65096, 65097, 65097, 65097, 65097, 65097, 65098, 65098, 65098, 65098, 65098, 65099, 65099, 65099, 65099, 65099, 65100, 65100, 65100, 65100, 65101, 65101, 65101, 65101, 65101, 65102, 65102, 65102, 65102, 65102, 65103, 65103, 65103, 65103, 65104, 65104, 65104, 65104, 65104, 65105, 65105, 65105, 65105, 65105, 65106, 65106, 65106, 65106, 65106, 65107, 65107, 65107, 65107, 65107, 65108, 65108, 65108, 65108, 65109, 65109, 65109, 65109, 65109, 65110, 65110, 65110, 65110, 65110, 65111, 65111, 65111, 65111, 65111, 65112, 65112, 65112, 65112, 65112, 65113, 65113, 65113, 65113, 65113, 65114, 65114, 65114, 65114, 65114, 65115, 65115, 65115, 65115, 65116, 65116, 65116, 65116, 65116, 65117, 65117, 65117, 65117, 65117, 65118, 65118, 65118, 65118, 65118, 65119, 65119, 65119, 65119, 65119, 65120, 65120, 65120, 65120, 65120, 65121, 65121, 65121, 65121, 65121, 65122, 65122, 65122, 65122, 65122, 65123, 65123, 65123, 65123, 65123, 65124, 65124, 65124, 65124, 65124, 65125, 65125, 65125, 65125, 65125, 65126, 65126, 65126, 65126, 65126, 65127, 65127, 65127, 65127, 65127, 65128, 65128, 65128, 65128, 65128, 65129, 65129, 65129, 65129, 65129, 65130, 65130, 65130, 65130, 65130, 65131, 65131, 65131, 65131, 65131, 65132, 65132, 65132, 65132, 65132, 65132, 65133, 65133, 65133, 65133, 65133, 65134, 65134, 65134, 65134, 65134, 65135, 65135, 65135, 65135, 65135, 65136, 65136, 65136, 65136, 65136, 65137, 65137, 65137, 65137, 65137, 65138, 65138, 65138, 65138, 65138, 65139, 65139, 65139, 65139, 65139, 65139, 65140, 65140, 65140, 65140, 65140, 65141, 65141, 65141, 65141, 65141, 65142, 65142, 65142, 65142, 65142, 65143, 65143, 65143, 65143, 65143, 65144, 65144, 65144, 65144, 65144, 65144, 65145, 65145, 65145, 65145, 65145, 65146, 65146, 65146, 65146, 65146, 65147, 65147, 65147, 65147, 65147, 65147, 65148, 65148, 65148, 65148, 65148, 65149, 65149, 65149, 65149, 65149, 65150, 65150, 65150, 65150, 65150, 65150, 65151, 65151, 65151, 65151, 65151, 65152, 65152, 65152, 65152, 65152, 65153, 65153, 65153, 65153, 65153, 65153, 65154, 65154, 65154, 65154, 65154, 65155, 65155, 65155, 65155, 65155, 65156, 65156, 65156, 65156, 65156, 65156, 65157, 65157, 65157, 65157, 65157, 65158, 65158, 65158, 65158, 65158, 65158, 65159, 65159, 65159, 65159, 65159, 65160, 65160, 65160, 65160, 65160, 65160, 65161, 65161, 65161, 65161, 65161, 65162, 65162, 65162, 65162, 65162, 65162, 65163, 65163, 65163, 65163, 65163, 65164, 65164, 65164, 65164, 65164, 65164, 65165, 65165, 65165, 65165, 65165, 65166, 65166, 65166, 65166, 65166, 65166, 65167, 65167, 65167, 65167, 65167, 65168, 65168, 65168, 65168, 65168, 65168, 65169, 65169, 65169, 65169, 65169, 65169, 65170, 65170, 65170, 65170, 65170, 65171, 65171, 65171, 65171, 65171, 65171, 65172, 65172, 65172, 65172, 65172, 65172, 65173, 65173, 65173, 65173, 65173, 65174, 65174, 65174, 65174, 65174, 65174, 65175, 65175, 65175, 65175, 65175, 65175, 65176, 65176, 65176, 65176, 65176, 65177, 65177, 65177, 65177, 65177, 65177, 65178, 65178, 65178, 65178, 65178, 65178, 65179, 65179, 65179, 65179, 65179, 65179, 65180, 65180, 65180, 65180, 65180, 65181, 65181, 65181, 65181, 65181, 65181, 65182, 65182, 65182, 65182, 65182, 65182, 65183, 65183, 65183, 65183, 65183, 65183, 65184, 65184, 65184, 65184, 65184, 65184, 65185, 65185, 65185, 65185, 65185, 65185, 65186, 65186, 65186, 65186, 65186, 65187, 65187, 65187, 65187, 65187, 65187, 65188, 65188, 65188, 65188, 65188, 65188, 65189, 65189, 65189, 65189, 65189, 65189, 65190, 65190, 65190, 65190, 65190, 65190, 65191, 65191, 65191, 65191, 65191, 65191, 65192, 65192, 65192, 65192, 65192, 65192, 65193, 65193, 65193, 65193, 65193, 65193, 65194, 65194, 65194, 65194, 65194, 65194, 65195, 65195, 65195, 65195, 65195, 65195, 65196, 65196, 65196, 65196, 65196, 65196, 65197, 65197, 65197, 65197, 65197, 65197, 65198, 65198, 65198, 65198, 65198, 65198, 65199, 65199, 65199, 65199, 65199, 65199, 65199, 65200, 65200, 65200, 65200, 65200, 65200, 65201, 65201, 65201, 65201, 65201, 65201, 65202, 65202, 65202, 65202, 65202, 65202, 65203, 65203, 65203, 65203, 65203, 65203, 65204, 65204, 65204, 65204, 65204, 65204, 65205, 65205, 65205, 65205, 65205, 65205, 65205, 65206, 65206, 65206, 65206, 65206, 65206, 65207, 65207, 65207, 65207, 65207, 65207, 65208, 65208, 65208, 65208, 65208, 65208, 65209, 65209, 65209, 65209, 65209, 65209, 65209, 65210, 65210, 65210, 65210, 65210, 65210, 65211, 65211, 65211, 65211, 65211, 65211, 65212, 65212, 65212, 65212, 65212, 65212, 65212, 65213, 65213, 65213, 65213, 65213, 65213, 65214, 65214, 65214, 65214, 65214, 65214, 65215, 65215, 65215, 65215, 65215, 65215, 65215, 65216, 65216, 65216, 65216, 65216, 65216, 65217, 65217, 65217, 65217, 65217, 65217, 65217, 65218, 65218, 65218, 65218, 65218, 65218, 65219, 65219, 65219, 65219, 65219, 65219, 65219, 65220, 65220, 65220, 65220, 65220, 65220, 65221, 65221, 65221, 65221, 65221, 65221, 65221, 65222, 65222, 65222, 65222, 65222, 65222, 65223, 65223, 65223, 65223, 65223, 65223, 65223, 65224, 65224, 65224, 65224, 65224, 65224, 65225, 65225, 65225, 65225, 65225, 65225, 65225, 65226, 65226, 65226, 65226, 65226, 65226, 65226, 65227, 65227, 65227, 65227, 65227, 65227, 65228, 65228, 65228, 65228, 65228, 65228, 65228, 65229, 65229, 65229, 65229, 65229, 65229, 65229, 65230, 65230, 65230, 65230, 65230, 65230, 65231, 65231, 65231, 65231, 65231, 65231, 65231, 65232, 65232, 65232, 65232, 65232, 65232, 65232, 65233, 65233, 65233, 65233, 65233, 65233, 65233, 65234, 65234, 65234, 65234, 65234, 65234, 65234, 65235, 65235, 65235, 65235, 65235, 65235, 65236, 65236, 65236, 65236, 65236, 65236, 65236, 65237, 65237, 65237, 65237, 65237, 65237, 65237, 65238, 65238, 65238, 65238, 65238, 65238, 65238, 65239, 65239, 65239, 65239, 65239, 65239, 65239, 65240, 65240, 65240, 65240, 65240, 65240, 65240, 65241, 65241, 65241, 65241, 65241, 65241, 65241, 65242, 65242, 65242, 65242, 65242, 65242, 65242, 65243, 65243, 65243, 65243, 65243, 65243, 65243, 65244, 65244, 65244, 65244, 65244, 65244, 65244, 65245, 65245, 65245, 65245, 65245, 65245, 65245, 65246, 65246, 65246, 65246, 65246, 65246, 65246, 65247, 65247, 65247, 65247, 65247, 65247, 65247, 65248, 65248, 65248, 65248, 65248, 65248, 65248, 65249, 65249, 65249, 65249, 65249, 65249, 65249, 65249, 65250, 65250, 65250, 65250, 65250, 65250, 65250, 65251, 65251, 65251, 65251, 65251, 65251, 65251, 65252, 65252, 65252, 65252, 65252, 65252, 65252, 65253, 65253, 65253, 65253, 65253, 65253, 65253, 65254, 65254, 65254, 65254, 65254, 65254, 65254, 65254, 65255, 65255, 65255, 65255, 65255, 65255, 65255, 65256, 65256, 65256, 65256, 65256, 65256, 65256, 65257, 65257, 65257, 65257, 65257, 65257, 65257, 65257, 65258, 65258, 65258, 65258, 65258, 65258, 65258, 65259, 65259, 65259, 65259, 65259, 65259, 65259, 65259, 65260, 65260, 65260, 65260, 65260, 65260, 65260, 65261, 65261, 65261, 65261, 65261, 65261, 65261, 65261, 65262, 65262, 65262, 65262, 65262, 65262, 65262, 65263, 65263, 65263, 65263, 65263, 65263, 65263, 65263, 65264, 65264, 65264, 65264, 65264, 65264, 65264, 65265, 65265, 65265, 65265, 65265, 65265, 65265, 65265, 65266, 65266, 65266, 65266, 65266, 65266, 65266, 65267, 65267, 65267, 65267, 65267, 65267, 65267, 65267, 65268, 65268, 65268, 65268, 65268, 65268, 65268, 65268, 65269, 65269, 65269, 65269, 65269, 65269, 65269, 65270, 65270, 65270, 65270, 65270, 65270, 65270, 65270, 65271, 65271, 65271, 65271, 65271, 65271, 65271, 65271, 65272, 65272, 65272, 65272, 65272, 65272, 65272, 65272, 65273, 65273, 65273, 65273, 65273, 65273, 65273, 65274, 65274, 65274, 65274, 65274, 65274, 65274, 65274, 65275, 65275, 65275, 65275, 65275, 65275, 65275, 65275, 65276, 65276, 65276, 65276, 65276, 65276, 65276, 65276, 65277, 65277, 65277, 65277, 65277, 65277, 65277, 65277, 65278, 65278, 65278, 65278, 65278, 65278, 65278, 65278, 65279, 65279, 65279, 65279, 65279, 65279, 65279, 65279, 65280, 65280, 65280, 65280, 65280, 65280, 65280, 65280, 65281, 65281, 65281, 65281, 65281, 65281, 65281, 65281, 65282, 65282, 65282, 65282, 65282, 65282, 65282, 65282, 65283, 65283, 65283, 65283, 65283, 65283, 65283, 65283, 65284, 65284, 65284, 65284, 65284, 65284, 65284, 65284, 65285, 65285, 65285, 65285, 65285, 65285, 65285, 65285, 65285, 65286, 65286, 65286, 65286, 65286, 65286, 65286, 65286, 65287, 65287, 65287, 65287, 65287, 65287, 65287, 65287, 65288, 65288, 65288, 65288, 65288, 65288, 65288, 65288, 65289, 65289, 65289, 65289, 65289, 65289, 65289, 65289, 65289, 65290, 65290, 65290, 65290, 65290, 65290, 65290, 65290, 65291, 65291, 65291, 65291, 65291, 65291, 65291, 65291, 65292, 65292, 65292, 65292, 65292, 65292, 65292, 65292, 65292, 65293, 65293, 65293, 65293, 65293, 65293, 65293, 65293, 65294, 65294, 65294, 65294, 65294, 65294, 65294, 65294, 65294, 65295, 65295, 65295, 65295, 65295, 65295, 65295, 65295, 65296, 65296, 65296, 65296, 65296, 65296, 65296, 65296, 65296, 65297, 65297, 65297, 65297, 65297, 65297, 65297, 65297, 65297, 65298, 65298, 65298, 65298, 65298, 65298, 65298, 65298, 65299, 65299, 65299, 65299, 65299, 65299, 65299, 65299, 65299, 65300, 65300, 65300, 65300, 65300, 65300, 65300, 65300, 65300, 65301, 65301, 65301, 65301, 65301, 65301, 65301, 65301, 65302, 65302, 65302, 65302, 65302, 65302, 65302, 65302, 65302, 65303, 65303, 65303, 65303, 65303, 65303, 65303, 65303, 65303, 65304, 65304, 65304, 65304, 65304, 65304, 65304, 65304, 65304, 65305, 65305, 65305, 65305, 65305, 65305, 65305, 65305, 65305, 65306, 65306, 65306, 65306, 65306, 65306, 65306, 65306, 65306, 65307, 65307, 65307, 65307, 65307, 65307, 65307, 65307, 65307, 65308, 65308, 65308, 65308, 65308, 65308, 65308, 65308, 65308, 65309, 65309, 65309, 65309, 65309, 65309, 65309, 65309, 65309, 65310, 65310, 65310, 65310, 65310, 65310, 65310, 65310, 65310, 65311, 65311, 65311, 65311, 65311, 65311, 65311, 65311, 65311, 65312, 65312, 65312, 65312, 65312, 65312, 65312, 65312, 65312, 65313, 65313, 65313, 65313, 65313, 65313, 65313, 65313, 65313, 65314, 65314, 65314, 65314, 65314, 65314, 65314, 65314, 65314, 65314, 65315, 65315, 65315, 65315, 65315, 65315, 65315, 65315, 65315, 65316, 65316, 65316, 65316, 65316, 65316, 65316, 65316, 65316, 65317, 65317, 65317, 65317, 65317, 65317, 65317, 65317, 65317, 65317, 65318, 65318, 65318, 65318, 65318, 65318, 65318, 65318, 65318, 65319, 65319, 65319, 65319, 65319, 65319, 65319, 65319, 65319, 65320, 65320, 65320, 65320, 65320, 65320, 65320, 65320, 65320, 65320, 65321, 65321, 65321, 65321, 65321, 65321, 65321, 65321, 65321, 65321, 65322, 65322, 65322, 65322, 65322, 65322, 65322, 65322, 65322, 65323, 65323, 65323, 65323, 65323, 65323, 65323, 65323, 65323, 65323, 65324, 65324, 65324, 65324, 65324, 65324, 65324, 65324, 65324, 65325, 65325, 65325, 65325, 65325, 65325, 65325, 65325, 65325, 65325, 65326, 65326, 65326, 65326, 65326, 65326, 65326, 65326, 65326, 65326, 65327, 65327, 65327, 65327, 65327, 65327, 65327, 65327, 65327, 65327, 65328, 65328, 65328, 65328, 65328, 65328, 65328, 65328, 65328, 65328, 65329, 65329, 65329, 65329, 65329, 65329, 65329, 65329, 65329, 65329, 65330, 65330, 65330, 65330, 65330, 65330, 65330, 65330, 65330, 65330, 65331, 65331, 65331, 65331, 65331, 65331, 65331, 65331, 65331, 65331, 65332, 65332, 65332, 65332, 65332, 65332, 65332, 65332, 65332, 65332, 65333, 65333, 65333, 65333, 65333, 65333, 65333, 65333, 65333, 65333, 65334, 65334, 65334, 65334, 65334, 65334, 65334, 65334, 65334, 65334, 65335, 65335, 65335, 65335, 65335, 65335, 65335, 65335, 65335, 65335, 65336, 65336, 65336, 65336, 65336, 65336, 65336, 65336, 65336, 65336, 65337, 65337, 65337, 65337, 65337, 65337, 65337, 65337, 65337, 65337, 65337, 65338, 65338, 65338, 65338, 65338, 65338, 65338, 65338, 65338, 65338, 65339, 65339, 65339, 65339, 65339, 65339, 65339, 65339, 65339, 65339, 65339, 65340, 65340, 65340, 65340, 65340, 65340, 65340, 65340, 65340, 65340, 65341, 65341, 65341, 65341, 65341, 65341, 65341, 65341, 65341, 65341, 65341, 65342, 65342, 65342, 65342, 65342, 65342, 65342, 65342, 65342, 65342, 65343, 65343, 65343, 65343, 65343, 65343, 65343, 65343, 65343, 65343, 65343, 65344, 65344, 65344, 65344, 65344, 65344, 65344, 65344, 65344, 65344, 65344, 65345, 65345, 65345, 65345, 65345, 65345, 65345, 65345, 65345, 65345, 65346, 65346, 65346, 65346, 65346, 65346, 65346, 65346, 65346, 65346, 65346, 65347, 65347, 65347, 65347, 65347, 65347, 65347, 65347, 65347, 65347, 65347, 65348, 65348, 65348, 65348, 65348, 65348, 65348, 65348, 65348, 65348, 65348, 65349, 65349, 65349, 65349, 65349, 65349, 65349, 65349, 65349, 65349, 65349, 65350, 65350, 65350, 65350, 65350, 65350, 65350, 65350, 65350, 65350, 65350, 65351, 65351, 65351, 65351, 65351, 65351, 65351, 65351, 65351, 65351, 65351, 65352, 65352, 65352, 65352, 65352, 65352, 65352, 65352, 65352, 65352, 65352, 65353, 65353, 65353, 65353, 65353, 65353, 65353, 65353, 65353, 65353, 65353, 65354, 65354, 65354, 65354, 65354, 65354, 65354, 65354, 65354, 65354, 65354, 65354, 65355, 65355, 65355, 65355, 65355, 65355, 65355, 65355, 65355, 65355, 65355, 65356, 65356, 65356, 65356, 65356, 65356, 65356, 65356, 65356, 65356, 65356, 65357, 65357, 65357, 65357, 65357, 65357, 65357, 65357, 65357, 65357, 65357, 65357, 65358, 65358, 65358, 65358, 65358, 65358, 65358, 65358, 65358, 65358, 65358, 65359, 65359, 65359, 65359, 65359, 65359, 65359, 65359, 65359, 65359, 65359, 65359, 65360, 65360, 65360, 65360, 65360, 65360, 65360, 65360, 65360, 65360, 65360, 65360, 65361, 65361, 65361, 65361, 65361, 65361, 65361, 65361, 65361, 65361, 65361, 65362, 65362, 65362, 65362, 65362, 65362, 65362, 65362, 65362, 65362, 65362, 65362, 65363, 65363, 65363, 65363, 65363, 65363, 65363, 65363, 65363, 65363, 65363, 65363, 65364, 65364, 65364, 65364, 65364, 65364, 65364, 65364, 65364, 65364, 65364, 65364, 65365, 65365, 65365, 65365, 65365, 65365, 65365, 65365, 65365, 65365, 65365, 65365, 65366, 65366, 65366, 65366, 65366, 65366, 65366, 65366, 65366, 65366, 65366, 65366, 65367, 65367, 65367, 65367, 65367, 65367, 65367, 65367, 65367, 65367, 65367, 65367, 65368, 65368, 65368, 65368, 65368, 65368, 65368, 65368, 65368, 65368, 65368, 65368, 65368, 65369, 65369, 65369, 65369, 65369, 65369, 65369, 65369, 65369, 65369, 65369, 65369, 65370, 65370, 65370, 65370, 65370, 65370, 65370, 65370, 65370, 65370, 65370, 65370, 65371, 65371, 65371, 65371, 65371, 65371, 65371, 65371, 65371, 65371, 65371, 65371, 65371, 65372, 65372, 65372, 65372, 65372, 65372, 65372, 65372, 65372, 65372, 65372, 65372, 65373, 65373, 65373, 65373, 65373, 65373, 65373, 65373, 65373, 65373, 65373, 65373, 65373, 65374, 65374, 65374, 65374, 65374, 65374, 65374, 65374, 65374, 65374, 65374, 65374, 65375, 65375, 65375, 65375, 65375, 65375, 65375, 65375, 65375, 65375, 65375, 65375, 65375, 65376, 65376, 65376, 65376, 65376, 65376, 65376, 65376, 65376, 65376, 65376, 65376, 65376, 65377, 65377, 65377, 65377, 65377, 65377, 65377, 65377, 65377, 65377, 65377, 65377, 65377, 65378, 65378, 65378, 65378, 65378, 65378, 65378, 65378, 65378, 65378, 65378, 65378, 65378, 65379, 65379, 65379, 65379, 65379, 65379, 65379, 65379, 65379, 65379, 65379, 65379, 65379, 65380, 65380, 65380, 65380, 65380, 65380, 65380, 65380, 65380, 65380, 65380, 65380, 65380, 65381, 65381, 65381, 65381, 65381, 65381, 65381, 65381, 65381, 65381, 65381, 65381, 65381, 65382, 65382, 65382, 65382, 65382, 65382, 65382, 65382, 65382, 65382, 65382, 65382, 65382, 65382, 65383, 65383, 65383, 65383, 65383, 65383, 65383, 65383, 65383, 65383, 65383, 65383, 65383, 65384, 65384, 65384, 65384, 65384, 65384, 65384, 65384, 65384, 65384, 65384, 65384, 65384, 65384, 65385, 65385, 65385, 65385, 65385, 65385, 65385, 65385, 65385, 65385, 65385, 65385, 65385, 65386, 65386, 65386, 65386, 65386, 65386, 65386, 65386, 65386, 65386, 65386, 65386, 65386, 65386, 65387, 65387, 65387, 65387, 65387, 65387, 65387, 65387, 65387, 65387, 65387, 65387, 65387, 65387, 65388, 65388, 65388, 65388, 65388, 65388, 65388, 65388, 65388, 65388, 65388, 65388, 65388, 65388, 65389, 65389, 65389, 65389, 65389, 65389, 65389, 65389, 65389, 65389, 65389, 65389, 65389, 65389, 65390, 65390, 65390, 65390, 65390, 65390, 65390, 65390, 65390, 65390, 65390, 65390, 65390, 65390, 65391, 65391, 65391, 65391, 65391, 65391, 65391, 65391, 65391, 65391, 65391, 65391, 65391, 65391, 65392, 65392, 65392, 65392, 65392, 65392, 65392, 65392, 65392, 65392, 65392, 65392, 65392, 65392, 65393, 65393, 65393, 65393, 65393, 65393, 65393, 65393, 65393, 65393, 65393, 65393, 65393, 65393, 65394, 65394, 65394, 65394, 65394, 65394, 65394, 65394, 65394, 65394, 65394, 65394, 65394, 65394, 65394, 65395, 65395, 65395, 65395, 65395, 65395, 65395, 65395, 65395, 65395, 65395, 65395, 65395, 65395, 65396, 65396, 65396, 65396, 65396, 65396, 65396, 65396, 65396, 65396, 65396, 65396, 65396, 65396, 65396, 65397, 65397, 65397, 65397, 65397, 65397, 65397, 65397, 65397, 65397, 65397, 65397, 65397, 65397, 65397, 65398, 65398, 65398, 65398, 65398, 65398, 65398, 65398, 65398, 65398, 65398, 65398, 65398, 65398, 65398, 65399, 65399, 65399, 65399, 65399, 65399, 65399, 65399, 65399, 65399, 65399, 65399, 65399, 65399, 65399, 65400, 65400, 65400, 65400, 65400, 65400, 65400, 65400, 65400, 65400, 65400, 65400, 65400, 65400, 65400, 65401, 65401, 65401, 65401, 65401, 65401, 65401, 65401, 65401, 65401, 65401, 65401, 65401, 65401, 65401, 65402, 65402, 65402, 65402, 65402, 65402, 65402, 65402, 65402, 65402, 65402, 65402, 65402, 65402, 65402, 65403, 65403, 65403, 65403, 65403, 65403, 65403, 65403, 65403, 65403, 65403, 65403, 65403, 65403, 65403, 65403, 65404, 65404, 65404, 65404, 65404, 65404, 65404, 65404, 65404, 65404, 65404, 65404, 65404, 65404, 65404, 65405, 65405, 65405, 65405, 65405, 65405, 65405, 65405, 65405, 65405, 65405, 65405, 65405, 65405, 65405, 65405, 65406, 65406, 65406, 65406, 65406, 65406, 65406, 65406, 65406, 65406, 65406, 65406, 65406, 65406, 65406, 65406, 65407, 65407, 65407, 65407, 65407, 65407, 65407, 65407, 65407, 65407, 65407, 65407, 65407, 65407, 65407, 65407, 65408, 65408, 65408, 65408, 65408, 65408, 65408, 65408, 65408, 65408, 65408, 65408, 65408, 65408, 65408, 65408, 65409, 65409, 65409, 65409, 65409, 65409, 65409, 65409, 65409, 65409, 65409, 65409, 65409, 65409, 65409, 65409, 65410, 65410, 65410, 65410, 65410, 65410, 65410, 65410, 65410, 65410, 65410, 65410, 65410, 65410, 65410, 65410, 65411, 65411, 65411, 65411, 65411, 65411, 65411, 65411, 65411, 65411, 65411, 65411, 65411, 65411, 65411, 65411, 65412, 65412, 65412, 65412, 65412, 65412, 65412, 65412, 65412, 65412, 65412, 65412, 65412, 65412, 65412, 65412, 65412, 65413, 65413, 65413, 65413, 65413, 65413, 65413, 65413, 65413, 65413, 65413, 65413, 65413, 65413, 65413, 65413, 65413, 65414, 65414, 65414, 65414, 65414, 65414, 65414, 65414, 65414, 65414, 65414, 65414, 65414, 65414, 65414, 65414, 65414, 65415, 65415, 65415, 65415, 65415, 65415, 65415, 65415, 65415, 65415, 65415, 65415, 65415, 65415, 65415, 65415, 65416, 65416, 65416, 65416, 65416, 65416, 65416, 65416, 65416, 65416, 65416, 65416, 65416, 65416, 65416, 65416, 65416, 65416, 65417, 65417, 65417, 65417, 65417, 65417, 65417, 65417, 65417, 65417, 65417, 65417, 65417, 65417, 65417, 65417, 65417, 65418, 65418, 65418, 65418, 65418, 65418, 65418, 65418, 65418, 65418, 65418, 65418, 65418, 65418, 65418, 65418, 65418, 65419, 65419, 65419, 65419, 65419, 65419, 65419, 65419, 65419, 65419, 65419, 65419, 65419, 65419, 65419, 65419, 65419, 65419, 65420, 65420, 65420, 65420, 65420, 65420, 65420, 65420, 65420, 65420, 65420, 65420, 65420, 65420, 65420, 65420, 65420, 65421, 65421, 65421, 65421, 65421, 65421, 65421, 65421, 65421, 65421, 65421, 65421, 65421, 65421, 65421, 65421, 65421, 65421, 65422, 65422, 65422, 65422, 65422, 65422, 65422, 65422, 65422, 65422, 65422, 65422, 65422, 65422, 65422, 65422, 65422, 65422, 65423, 65423, 65423, 65423, 65423, 65423, 65423, 65423, 65423, 65423, 65423, 65423, 65423, 65423, 65423, 65423, 65423, 65423, 65424, 65424, 65424, 65424, 65424, 65424, 65424, 65424, 65424, 65424, 65424, 65424, 65424, 65424, 65424, 65424, 65424, 65424, 65424, 65425, 65425, 65425, 65425, 65425, 65425, 65425, 65425, 65425, 65425, 65425, 65425, 65425, 65425, 65425, 65425, 65425, 65425, 65426, 65426, 65426, 65426, 65426, 65426, 65426, 65426, 65426, 65426, 65426, 65426, 65426, 65426, 65426, 65426, 65426, 65426, 65426, 65427, 65427, 65427, 65427, 65427, 65427, 65427, 65427, 65427, 65427, 65427, 65427, 65427, 65427, 65427, 65427, 65427, 65427, 65427, 65428, 65428, 65428, 65428, 65428, 65428, 65428, 65428, 65428, 65428, 65428, 65428, 65428, 65428, 65428, 65428, 65428, 65428, 65428, 65429, 65429, 65429, 65429, 65429, 65429, 65429, 65429, 65429, 65429, 65429, 65429, 65429, 65429, 65429, 65429, 65429, 65429, 65429, 65430, 65430, 65430, 65430, 65430, 65430, 65430, 65430, 65430, 65430, 65430, 65430, 65430, 65430, 65430, 65430, 65430, 65430, 65430, 65431, 65431, 65431, 65431, 65431, 65431, 65431, 65431, 65431, 65431, 65431, 65431, 65431, 65431, 65431, 65431, 65431, 65431, 65431, 65431, 65432, 65432, 65432, 65432, 65432, 65432, 65432, 65432, 65432, 65432, 65432, 65432, 65432, 65432, 65432, 65432, 65432, 65432, 65432, 65433, 65433, 65433, 65433, 65433, 65433, 65433, 65433, 65433, 65433, 65433, 65433, 65433, 65433, 65433, 65433, 65433, 65433, 65433, 65433, 65434, 65434, 65434, 65434, 65434, 65434, 65434, 65434, 65434, 65434, 65434, 65434, 65434, 65434, 65434, 65434, 65434, 65434, 65434, 65434, 65435, 65435, 65435, 65435, 65435, 65435, 65435, 65435, 65435, 65435, 65435, 65435, 65435, 65435, 65435, 65435, 65435, 65435, 65435, 65435, 65435, 65436, 65436, 65436, 65436, 65436, 65436, 65436, 65436, 65436, 65436, 65436, 65436, 65436, 65436, 65436, 65436, 65436, 65436, 65436, 65436, 65437, 65437, 65437, 65437, 65437, 65437, 65437, 65437, 65437, 65437, 65437, 65437, 65437, 65437, 65437, 65437, 65437, 65437, 65437, 65437, 65437, 65438, 65438, 65438, 65438, 65438, 65438, 65438, 65438, 65438, 65438, 65438, 65438, 65438, 65438, 65438, 65438, 65438, 65438, 65438, 65438, 65438, 65439, 65439, 65439, 65439, 65439, 65439, 65439, 65439, 65439, 65439, 65439, 65439, 65439, 65439, 65439, 65439, 65439, 65439, 65439, 65439, 65439, 65440, 65440, 65440, 65440, 65440, 65440, 65440, 65440, 65440, 65440, 65440, 65440, 65440, 65440, 65440, 65440, 65440, 65440, 65440, 65440, 65440, 65441, 65441, 65441, 65441, 65441, 65441, 65441, 65441, 65441, 65441, 65441, 65441, 65441, 65441, 65441, 65441, 65441, 65441, 65441, 65441, 65441, 65441, 65442, 65442, 65442, 65442, 65442, 65442, 65442, 65442, 65442, 65442, 65442, 65442, 65442, 65442, 65442, 65442, 65442, 65442, 65442, 65442, 65442, 65442, 65443, 65443, 65443, 65443, 65443, 65443, 65443, 65443, 65443, 65443, 65443, 65443, 65443, 65443, 65443, 65443, 65443, 65443, 65443, 65443, 65443, 65443, 65444, 65444, 65444, 65444, 65444, 65444, 65444, 65444, 65444, 65444, 65444, 65444, 65444, 65444, 65444, 65444, 65444, 65444, 65444, 65444, 65444, 65444, 65445, 65445, 65445, 65445, 65445, 65445, 65445, 65445, 65445, 65445, 65445, 65445, 65445, 65445, 65445, 65445, 65445, 65445, 65445, 65445, 65445, 65445, 65445, 65446, 65446, 65446, 65446, 65446, 65446, 65446, 65446, 65446, 65446, 65446, 65446, 65446, 65446, 65446, 65446, 65446, 65446, 65446, 65446, 65446, 65446, 65446, 65447, 65447, 65447, 65447, 65447, 65447, 65447, 65447, 65447, 65447, 65447, 65447, 65447, 65447, 65447, 65447, 65447, 65447, 65447, 65447, 65447, 65447, 65447, 65448, 65448, 65448, 65448, 65448, 65448, 65448, 65448, 65448, 65448, 65448, 65448, 65448, 65448, 65448, 65448, 65448, 65448, 65448, 65448, 65448, 65448, 65448, 65449, 65449, 65449, 65449, 65449, 65449, 65449, 65449, 65449, 65449, 65449, 65449, 65449, 65449, 65449, 65449, 65449, 65449, 65449, 65449, 65449, 65449, 65449, 65450, 65450, 65450, 65450, 65450, 65450, 65450, 65450, 65450, 65450, 65450, 65450, 65450, 65450, 65450, 65450, 65450, 65450, 65450, 65450, 65450, 65450, 65450, 65450, 65451, 65451, 65451, 65451, 65451, 65451, 65451, 65451, 65451, 65451, 65451, 65451, 65451, 65451, 65451, 65451, 65451, 65451, 65451, 65451, 65451, 65451, 65451, 65451, 65452, 65452, 65452, 65452, 65452, 65452, 65452, 65452, 65452, 65452, 65452, 65452, 65452, 65452, 65452, 65452, 65452, 65452, 65452, 65452, 65452, 65452, 65452, 65452, 65452, 65453, 65453, 65453, 65453, 65453, 65453, 65453, 65453, 65453, 65453, 65453, 65453, 65453, 65453, 65453, 65453, 65453, 65453, 65453, 65453, 65453, 65453, 65453, 65453, 65453, 65454, 65454, 65454, 65454, 65454, 65454, 65454, 65454, 65454, 65454, 65454, 65454, 65454, 65454, 65454, 65454, 65454, 65454, 65454, 65454, 65454, 65454, 65454, 65454, 65454, 65455, 65455, 65455, 65455, 65455, 65455, 65455, 65455, 65455, 65455, 65455, 65455, 65455, 65455, 65455, 65455, 65455, 65455, 65455, 65455, 65455, 65455, 65455, 65455, 65455, 65456, 65456, 65456, 65456, 65456, 65456, 65456, 65456, 65456, 65456, 65456, 65456, 65456, 65456, 65456, 65456, 65456, 65456, 65456, 65456, 65456, 65456, 65456, 65456, 65456, 65456, 65457, 65457, 65457, 65457, 65457, 65457, 65457, 65457, 65457, 65457, 65457, 65457, 65457, 65457, 65457, 65457, 65457, 65457, 65457, 65457, 65457, 65457, 65457, 65457, 65457, 65458, 65458, 65458, 65458, 65458, 65458, 65458, 65458, 65458, 65458, 65458, 65458, 65458, 65458, 65458, 65458, 65458, 65458, 65458, 65458, 65458, 65458, 65458, 65458, 65458, 65458, 65458, 65459, 65459, 65459, 65459, 65459, 65459, 65459, 65459, 65459, 65459, 65459, 65459, 65459, 65459, 65459, 65459, 65459, 65459, 65459, 65459, 65459, 65459, 65459, 65459, 65459, 65459, 65460, 65460, 65460, 65460, 65460, 65460, 65460, 65460, 65460, 65460, 65460, 65460, 65460, 65460, 65460, 65460, 65460, 65460, 65460, 65460, 65460, 65460, 65460, 65460, 65460, 65460, 65460, 65461, 65461, 65461, 65461, 65461, 65461, 65461, 65461, 65461, 65461, 65461, 65461, 65461, 65461, 65461, 65461, 65461, 65461, 65461, 65461, 65461, 65461, 65461, 65461, 65461, 65461, 65461, 65461, 65462, 65462, 65462, 65462, 65462, 65462, 65462, 65462, 65462, 65462, 65462, 65462, 65462, 65462, 65462, 65462, 65462, 65462, 65462, 65462, 65462, 65462, 65462, 65462, 65462, 65462, 65462, 65463, 65463, 65463, 65463, 65463, 65463, 65463, 65463, 65463, 65463, 65463, 65463, 65463, 65463, 65463, 65463, 65463, 65463, 65463, 65463, 65463, 65463, 65463, 65463, 65463, 65463, 65463, 65463, 65464, 65464, 65464, 65464, 65464, 65464, 65464, 65464, 65464, 65464, 65464, 65464, 65464, 65464, 65464, 65464, 65464, 65464, 65464, 65464, 65464, 65464, 65464, 65464, 65464, 65464, 65464, 65464, 65464, 65465, 65465, 65465, 65465, 65465, 65465, 65465, 65465, 65465, 65465, 65465, 65465, 65465, 65465, 65465, 65465, 65465, 65465, 65465, 65465, 65465, 65465, 65465, 65465, 65465, 65465, 65465, 65465, 65465, 65466, 65466, 65466, 65466, 65466, 65466, 65466, 65466, 65466, 65466, 65466, 65466, 65466, 65466, 65466, 65466, 65466, 65466, 65466, 65466, 65466, 65466, 65466, 65466, 65466, 65466, 65466, 65466, 65466, 65467, 65467, 65467, 65467, 65467, 65467, 65467, 65467, 65467, 65467, 65467, 65467, 65467, 65467, 65467, 65467, 65467, 65467, 65467, 65467, 65467, 65467, 65467, 65467, 65467, 65467, 65467, 65467, 65467, 65467, 65468, 65468, 65468, 65468, 65468, 65468, 65468, 65468, 65468, 65468, 65468, 65468, 65468, 65468, 65468, 65468, 65468, 65468, 65468, 65468, 65468, 65468, 65468, 65468, 65468, 65468, 65468, 65468, 65468, 65468, 65469, 65469, 65469, 65469, 65469, 65469, 65469, 65469, 65469, 65469, 65469, 65469, 65469, 65469, 65469, 65469, 65469, 65469, 65469, 65469, 65469, 65469, 65469, 65469, 65469, 65469, 65469, 65469, 65469, 65469, 65469, 65470, 65470, 65470, 65470, 65470, 65470, 65470, 65470, 65470, 65470, 65470, 65470, 65470, 65470, 65470, 65470, 65470, 65470, 65470, 65470, 65470, 65470, 65470, 65470, 65470, 65470, 65470, 65470, 65470, 65470, 65470, 65471, 65471, 65471, 65471, 65471, 65471, 65471, 65471, 65471, 65471, 65471, 65471, 65471, 65471, 65471, 65471, 65471, 65471, 65471, 65471, 65471, 65471, 65471, 65471, 65471, 65471, 65471, 65471, 65471, 65471, 65471, 65472, 65472, 65472, 65472, 65472, 65472, 65472, 65472, 65472, 65472, 65472, 65472, 65472, 65472, 65472, 65472, 65472, 65472, 65472, 65472, 65472, 65472, 65472, 65472, 65472, 65472, 65472, 65472, 65472, 65472, 65472, 65472, 65473, 65473, 65473, 65473, 65473, 65473, 65473, 65473, 65473, 65473, 65473, 65473, 65473, 65473, 65473, 65473, 65473, 65473, 65473, 65473, 65473, 65473, 65473, 65473, 65473, 65473, 65473, 65473, 65473, 65473, 65473, 65473, 65473, 65474, 65474, 65474, 65474, 65474, 65474, 65474, 65474, 65474, 65474, 65474, 65474, 65474, 65474, 65474, 65474, 65474, 65474, 65474, 65474, 65474, 65474, 65474, 65474, 65474, 65474, 65474, 65474, 65474, 65474, 65474, 65474, 65474, 65475, 65475, 65475, 65475, 65475, 65475, 65475, 65475, 65475, 65475, 65475, 65475, 65475, 65475, 65475, 65475, 65475, 65475, 65475, 65475, 65475, 65475, 65475, 65475, 65475, 65475, 65475, 65475, 65475, 65475, 65475, 65475, 65475, 65476, 65476, 65476, 65476, 65476, 65476, 65476, 65476, 65476, 65476, 65476, 65476, 65476, 65476, 65476, 65476, 65476, 65476, 65476, 65476, 65476, 65476, 65476, 65476, 65476, 65476, 65476, 65476, 65476, 65476, 65476, 65476, 65476, 65476, 65476, 65477, 65477, 65477, 65477, 65477, 65477, 65477, 65477, 65477, 65477, 65477, 65477, 65477, 65477, 65477, 65477, 65477, 65477, 65477, 65477, 65477, 65477, 65477, 65477, 65477, 65477, 65477, 65477, 65477, 65477, 65477, 65477, 65477, 65477, 65478, 65478, 65478, 65478, 65478, 65478, 65478, 65478, 65478, 65478, 65478, 65478, 65478, 65478, 65478, 65478, 65478, 65478, 65478, 65478, 65478, 65478, 65478, 65478, 65478, 65478, 65478, 65478, 65478, 65478, 65478, 65478, 65478, 65478, 65478, 65478, 65479, 65479, 65479, 65479, 65479, 65479, 65479, 65479, 65479, 65479, 65479, 65479, 65479, 65479, 65479, 65479, 65479, 65479, 65479, 65479, 65479, 65479, 65479, 65479, 65479, 65479, 65479, 65479, 65479, 65479, 65479, 65479, 65479, 65479, 65479, 65479, 65480, 65480, 65480, 65480, 65480, 65480, 65480, 65480, 65480, 65480, 65480, 65480, 65480, 65480, 65480, 65480, 65480, 65480, 65480, 65480, 65480, 65480, 65480, 65480, 65480, 65480, 65480, 65480, 65480, 65480, 65480, 65480, 65480, 65480, 65480, 65480, 65481, 65481, 65481, 65481, 65481, 65481, 65481, 65481, 65481, 65481, 65481, 65481, 65481, 65481, 65481, 65481, 65481, 65481, 65481, 65481, 65481, 65481, 65481, 65481, 65481, 65481, 65481, 65481, 65481, 65481, 65481, 65481, 65481, 65481, 65481, 65481, 65481, 65481, 65482, 65482, 65482, 65482, 65482, 65482, 65482, 65482, 65482, 65482, 65482, 65482, 65482, 65482, 65482, 65482, 65482, 65482, 65482, 65482, 65482, 65482, 65482, 65482, 65482, 65482, 65482, 65482, 65482, 65482, 65482, 65482, 65482, 65482, 65482, 65482, 65482, 65483, 65483, 65483, 65483, 65483, 65483, 65483, 65483, 65483, 65483, 65483, 65483, 65483, 65483, 65483, 65483, 65483, 65483, 65483, 65483, 65483, 65483, 65483, 65483, 65483, 65483, 65483, 65483, 65483, 65483, 65483, 65483, 65483, 65483, 65483, 65483, 65483, 65483, 65483, 65484, 65484, 65484, 65484, 65484, 65484, 65484, 65484, 65484, 65484, 65484, 65484, 65484, 65484, 65484, 65484, 65484, 65484, 65484, 65484, 65484, 65484, 65484, 65484, 65484, 65484, 65484, 65484, 65484, 65484, 65484, 65484, 65484, 65484, 65484, 65484, 65484, 65484, 65484, 65484, 65485, 65485, 65485, 65485, 65485, 65485, 65485, 65485, 65485, 65485, 65485, 65485, 65485, 65485, 65485, 65485, 65485, 65485, 65485, 65485, 65485, 65485, 65485, 65485, 65485, 65485, 65485, 65485, 65485, 65485, 65485, 65485, 65485, 65485, 65485, 65485, 65485, 65485, 65485, 65485, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65486, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65487, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65488, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65489, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65490, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65491, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65492, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65493, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65494, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65495, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65496, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65497, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65498, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65499, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65500, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65501, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65502, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65503, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65504, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65505, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65506, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65507, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65508, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65509, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65510, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65511, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65512, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65513, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65514, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65515, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65516, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65517, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65518, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65519, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65520, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65521, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65522, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65523, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65524, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65525, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65526, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65527, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65528, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65529, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65530, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65531, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65532, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65533, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65534, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65535, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536, 65536);
end Sigmoid_Package;